`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
OMrdsrRpEttWODluC0AG3g/S5UKDr70bMwdgbqGF2RcL3xQFKYSyWp8fy2bHCB0EwAyCuxzOK/Q4
6r+SZfIUdA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
k2s7EWMhwIf9qGlEYH6Z9DmMZaK4vgWvIZZQxDcKCuHnkjHbD4/U7j76EMOamepLlmmJnKhUAdRO
dc+uAzJqa3NzMdAPJFre2fJTMQMEWzu/4dgityBiSUTOj+K+5pEFBnHCWSnQ5UzqFIY1yOb2/YZD
IG6YTCJbciIYaWhqK9s=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aILjgC2GmUyiU4AsUQ07DWXQjEHi3V5qONJrWxkXz62EwqxUiX7OkROoeH9DhNSRuL+w/JovcdHp
AnOkZd9mV20DGVARKPB0eQfKRK0AWUhYPWUtiiWeRu8Z+7BUxCklK5emK5hmSewVxkSJFo0so5mo
/3ixidv16V3WOQkjFJ0=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
f+rdl3qbw8Vh2sCsDZzrVbRhJv2vRjOjuOu9zad0VWeE/e0Kmt5X3+pZuwP1ihdaCNr0JAv3T12B
BeKSWuge5Jn1lRRnMDmqWo3VK/WtHWjPLg77Ld95Cw/UnVXF1nR8KwOwf1TsfRJJ90g2LFlsFCsO
htIB5UnYmtD/jtJQ7rqrR0vF5Ld08rcqInLs3GGqZDfE0y6HY1xbFDFdv2mHJmwV2wNo5H6ajr92
oLgFQJdGC14cOlecPHiyWr5oN06TlRrVu09xv57BRAuANqqr01cY4Hi1738LtV5zMIVnYvAgn7C1
n2jLIBA/dB+md2J//8MNc6k4rbbYTPpAbsJtvg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HIRSbdFYfaAF5GWQP4bTR1MpBjfvtA2Z+pbC6p3lNvvLlskzokTZ36tImVNUOW1pfCk899YaeKwq
TTiJDjb4JbOTrC9mCN1hx8O6tnLsEAYOGznzptkEtOSTHT9CyvXvtK11ZA5BmUsjolGm8yaYHIEo
UOS5B+SJRFWTGrho8hQ1WIDzGNytXdeuN+o4EUgHODMSlLFJSNdTZ0ne2PNM0dHMuiaGZQ9fsQo+
Y37J7Y+G9kPvZqUMJ9UyOGHZKySEPKY01qYx50ZsDjRXMKAI+B9AxUEB0IAl23nhNntbxobSir3F
rxd22+M0inY3utkXvyZJIFPfywY8ztrZOCDPlw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ltl0Tbg4fzfpcs5GkvjMeLedXpUr19ejb9G7kWMD8rRS1iPgypVcWiB2sDOnc2uWRfwgbvUtcLc6
QKoNQ7c7VYrt28FZQhVBJuhX8D6ipRuXrRhdRnNcY4d2SovB/6tZxv2U9LOTtPhivmr5egDbBE6Y
E3IkK7PsH1klzQySamoislPGqjg/NSgSWMDtjcSofaE7bKNbmUozSGqkROvv4uMmWcGd0wXrSd/1
YYlP/rPsSMe+OTsGDGElMp3uovABUt2G5v2eUUr586WGPnynPC4UYifriLnU7cAuyNfM/OI+oOe4
BBF66x/+pBsG0h2FnbXpUvNTUnqAl+APQ8CA7Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 261312)
`protect data_block
bIaiZoda0TAY/6wbCHXe/1MAWEWNwgC+5l8nn0EGf9cqAMAX3YeuDqPy7WAXNv/bcIaW+RliSc3k
ls6lQ3+8Q7VPPCcHWr6VMJ+q1u/JssFrX8zwN2mN/kx+8f8W8thrDRNljqzhUbOSRqMGKo2t29Pz
TJGWvRWzkm3OTHHFCV2fobtnOH10b19hB7sQBOeSfrhEVPLE+8oi0ThwpR/NR0IQCN6McMW6MHRb
Au7F5kQyuXGeZL2MwUSnGZFV5OyocyaFm/2xxbK4BCXVcPIKxJ13/rtgqnjEZBz/rzR5V/WS08fb
PgjYtwW3h5DhLMa6Uqajul0NVoQCNMkORKDUaEZ8deE1Zth75IEmjwBNdZFFhjQeYLyCsQ435jbC
KQ5qIAQAPcMaMeFA9c2EY4Yqm/zK2AWJLTdOcpUFkVFxjC04q9Yt1k3Qt7nOWJOkBihX8vrnVuap
I1VRgYygFNlIheu6IyFf8N3Nq/GiMSe9OsUjhZMFb05QqK+oeXg0nhdpJBZChY3M9u5QEv3pooU0
dQ8XHXpV/gSh/iee1voNcKwl6z7KgPFQyzUeRHEzzsa28jgGlpZCxrPpTctHlwQMl32vwb+UIRua
+KohSB3PDRea3znX3Iytm7oO7RO+fVCP4qpQVcyDVxVvsiUd2u01Dx5mdvSmN47g4mjzE6aGIzhg
E6vdu4S6eKswXdEaDQk2w7Z8uP+CYyKWKQOr4eGiIwVgFxBEIYirflhnfCelSoCBz9X600YEDq7X
n/u7V982jAUbTO/LyImO+LUpK1m8q4Cr0kHRZ0gDriACpDbxrWcvwlFWo8X3L2UiHN0aHjlXv7xU
6mHRA0ZqvcVkPxQjGmNV6+elX19vWDGv971znZ0YGz0VHOE30Tnv1TKhFWkW38dUfYOGO2YvRHC+
ysIVY/cuNzU1r4+LuWjHg9mdw9Ax9BDyLYknzLub+RbjuqFKg9cPbR3S5dwYk1N6g1ZPSQauGEwz
IxMvK2i7zKCdFcA+BrkMibO4jbB3dQ3Z2QfZdtTaLbUrEfGj7LMFH46+g4hi/uLbzvg+xYpp3g8h
7gXqX9hlWl6i88w9KeS46KFPKnQ0dR86KVKrJWa7IOHbDKeSqiqSQGPIEExNyKneTDZsW+lc5Wkh
qHtuvXO7bWEzZOWUzpYe61Ep36oUZXXvW0JBhGXvNE7ZItQkHuBV+oEQBYaLcm2jOwHc5TXRPjQd
PcKTcUqBOYdmC4ElNgoH6cqhzQV4nGnO7yweGxxRwgwtltipLonp7zaFhC0Eppb6JJ60pWRcjiU4
wUehzb6I8gtzEVLX+QgZdSjX9PtHDrN/Ljn39ihb1VorHPBLPqOeF0EwJ+M6s0kMppSSfMgt+5wS
7CYCvvBGPOcxUcXEA6n5Y+2t11QYpUMMmTpgfnSJOlW09DROuMMVNn2LIsSuUjydh1ihJfRFUmmD
2XpsVUJpXUH8yizMeh4nuKbVbgaFwQJm2toRZ0rpEXyjuVMAzYRLS/JWwlaSeUc+BId36O1dunHl
dfCaOx8s5luWVI21wGTzAZvcF2D0w1EtUFg9J/Q62POFVmy71IYFH4A0qXY4ZXOmD8NUq2bxWZVr
NnD1Ma5XrJ/oXs03uwnBqZ3I26V/hFKbDl476gdpUxr+oQgDPzo+1raCNYXRtG8EKeLeUUuQkmqk
AtF+Je0Yyn1Y62VleaC2sZReRLazVZT0/dkq46homQl9s5xSv9H3T9fa7+Wu5GuW80EiQfW6RqoB
Lu5wbIfvtIDrXvMEkj4pl3yvdNyrcC84MC3aWonK7G2CZEuLsDbZPFAg1Jt3o2hdwhYKU5CV/kqm
8rNK8PamCF3H3Sru9vt07Cmyl6OuIiytOSbir8zKRldVZ5p83Soqpc5/vwa+PPBR8oaGMKLiQ7xA
/M8/I5qb+pNxSteMeUWzBIEYR6Yfj9ANM7iGVQeh+PiqDk2Q8CwfHnvirszpanp2HkxA2p2+2t+n
AfFzPHmmmMRxogPC85UXksKCg2shY81Z5pLluxWcqQwm9FCf/yVd6sgFFh1AQc91uzJa1oClbSS3
NuFTWAb2u4RiFfdMhowFzCc8KVsxkvhvRfe9/XL7eUNAF03w/2hlwCrc3eI/oCT+fApvJ75/lg70
3RXbvgCq3i33KLkXNN+XHEqf1WVLGMYINQlsx2TdnCY+0AaLe1xoiTOY5J0NnBkrNEAzYT8YGE2T
vsjf9MhGmObeL8WkiaZwlvKjTbV6EjfDsf6mz9YFEW/HTrns3WA9FRbzENbbt+AaUvq1E3bksTO+
d1OkmzzGj82KZ3Jam9JcwuBOXGbZb9DeaV9ZcHjW3MiCu76u90JWtmc6vFjySJkUamEMqG4eOzvq
XYZtnQmo6iwTKV+XIzu2Cjd+BOrnM/rDjk9YK4ldLGsJc7fCXmiUH1pvMaPLxrbZX8c1SFn6wpjY
kQVCZSyl9uGmtm6/MAaS7Gcfhqpc1zIHLmS+MzAUPzK2ULFAr2F87g1ImhQWT3X4dVQY5blhrw74
W6IIH8ZYwGk2EFGmln4YlEdZYB67nPIHl1Ua5ziU1llQs0sqn+VCeBI5aCtvT1ZLygdMGGMOCFpT
eSkSRwnsXoWNyTTMJbFF9cArT9uo31L3ZU3qSj+OWInLjRlFkSUxlK41+DXG4g7MEj64pKjTxysp
ihUGg8TgcHoNkENsl48fmIgFtVPS3FoYEtfc615bIERQ2ogS0o8KkibuY6oBq/vSVY/K+MLzuTbd
qGZ6chEm9nq4FDAavigv+zG7y2d4BErDbBmFYYPbIp7nMDCvEMl5/7MFLtol6CZPiNFGYumuR/0m
ePT4Pua+29L6kO5RkZY4kSMIRcAX2XZcAdCUUGRs+lKTk+ZWD2EEFA7iO9dr9TAsyE0jMVeJ98e+
3WqVnzan6WmDKw+QuisJjb+N2bRahELkmIgl0TcYkO2QVf8jADnUJbWxYKd+yaIkisu5fe7e2MXN
v/B6CGqoyf69Bdy+5fsNHIYgBajOHSTflS8uBkkdygcp8DU5+m36tgQfzZKEROw5D/ExAX9Gyo8B
YYi2EdceZm+o4gDfYxh/wjpHU0D1YHAlrnTSpsbCYbRdwQlbLbKRVMlyBQcG63rMU72PEz+nzcNb
/0v6QL2M+GeJi2+LQe3rZV+gwPnSQVGJXZfJ6yxyTidTjYwLUW60Gzs2h8mJQynGsmIGIfn/bTNi
EY75JqO5Cua5qcmmCF+01Caj9p3YlQxJ3tmPJhxkTzcADwM5BdOtbsWK7ZtQ65c7b/UYKsMoRgEz
N6CDEOu1HYKAasJn6rmTu/itjHcqbpdWRKp9/jmO0xxt/WaW2ETp0dPf3atgvFeLhh9Z65T0q82H
DQpY47VamTLVlmfB1PRlTLUu1iTZWw3mqHJ3ijLzxBDUSbapmKkLU0MW01192ZcAvI3MJCK4Aj+K
gdeESkba70T5Zbv4k6fH8OWR0t6hnjyemYJO1yweEPzq9jRpca2o61SRfs1W/JG0y9nwBZKSRvJN
avLI55eNfsXxwtpA8jaNs4Ozjns1/cvO2PxcMyqyyygzhs5/Zn93qGQXNFSDoNaAXyy2cXcsPlKc
2L1wpNgitahrZLZVB762Rh8+JQktv3riM4O4kW5Fr5m3QOQTdT05eR1QoMhUCiIP4a4uYEbjv1Ua
igGaqTm+RwqjsUuReXkuItv4nsfeEgYAtDtlVFtLssVeqpvKF8loTvEweVl9+zSMwjbIxP5K+Y0m
H+ZjbQMYoFicR4TNh3yKet0XF10jXBIm/NO0JX5vtFOFrbIP+XEbAFTcrmIOOvrYOuHK0bBk01EJ
lUa2cASC5g+BchHHJqz+XRr65fTAYq1ZaiuZT5lgmF488P5E0fRd8UOr7+QSs+3Kzj40bjP9OM9n
JK6IwwnlFVjHCSJnJp0j4lj1uFWCcCiM9ElH8qpMjl0vTGN32ZPsC/ws8nSoDPLXn8nTaMcglWmK
77wsME3MfDJJQ/vfGNcg8zvafwm0WBYX4RiSm9a74oG4kMsbcGMluHU/Cw3crpjmmIXQ1mKSsHne
ZEpRRx8PL/bWyaSFuhxB4F85+VeFS1YM48YZUgq77e0i4SYs/cRfH4HqloLiN3EgdljWej2qth7/
3tKc5HzcmtGa2azZTY710tuz6/XCprN3CW3hC/n2xT8bpbzTr0Y/DLtxttSeZ+7KmarEm3prMud8
SZCU2HNtEZv+5jBR2iVk3JqIk5TMq70uxASAX6WHb7NYxFUmmk7HGWUt+4JZyYZn1mrvNw9YgNXn
KGN0nq07tOrbTkunJ9mUp7atRsKdBug0acw+7E3Uh9s+TENUZFiHD7nRj1Cx/cCFOBYq+wbqDWfz
zoefHXcVnednhVJ0qSx960XB3p+ddPyKnAd7hFgF1Y9bhwazlxekFi9jQl30kJFt6IlUebOkzCU1
qfDWIOfLR+o2K2FwnmwTj9AQekjFzA1O/fK0xF/XvbDmn8BzQSD+C6gd4Hqs/2ldaHd9e5Cvm3el
1I0IR7aeVEJaF1niFB4iWnH/0lAvZXIlbuY+eTdPO5sbkDIVbvhKllrc5OMAdqGPhGh+XoVVS4Go
Wxm62uv547U9ToUrYUgU3ii1DjpjGHb9b7SExiIOiTUYkUG8GKBidl95+5w+OvX1n2WEz7ZqLaS6
lk+eSPnrApigSUrwltUqmZgKjUXGUK5oy5dVLl/3UHew5wAe2SWf17AaolQdysp42rz1E1O6hru2
KMhIkaEqrn1z4vagsRvuUzI25LuaDFxkOqs9sebFz1KIFBRG/tihFSxhTvEZN2oXmVVe30qN/fdy
d3tMdpvoWsB5FyqdZMIDpRxlLqZuDtK+lPxM/8eatdw/jLeX3NYwCNrBBmYL5YC6kpnkALAHYypG
A6MZZB2n/xl53JBPOHN2P3Ej+NE1K5fum0DA5yh8vFZ41piynRhUNDpUmhPmHqWw9gGbiYPDAyVh
eV5yXc0+Ot8AQADp/t0cjPQumTZpu1G3ooaDDCXKHsLBSfKMtIYpAV7ddX+OTt/AEds4PvWuBeYc
B1EwZzdLQxFRPlWsH23oUdXvVVYzU5kLAkW6CYLMH1zLWMw1+baW8B0ok4FMlGKjAqwGnfg5opo1
O3+Jmy0UZCP5xDZHNsnJ5fDCm8gsyjJCfS+ILZCf+f7EUx+gNyT6pqFteeIofnWhwzBhVcFOVMly
+FNZYX5DXhLOMl0zWLbYVA1JYpD35rmgVzYEPWDkFxgsxdMLO+vsEIX7A+epocDQoUXcvxabxT/c
ZrAG111so3fFWFovu+HkrSKTdjt75i+31w3VNZJ69JXZ/Hr3hgHr03VCKljdk7UL+gzB+NG0huEH
0RF4H1At7/oGsGKgZcyh5w70QrxlyT/3ETnVXPjdd4BiPaPG9/MjbbtsMObQCWF1HJ9SDRhq1P4a
JRKnMuNaHD1k4EJj6c0I+TZFcF1kSaex7GI2CFMnfvOD5ax9LDIitRtmg9ywuvttPcynR9kPpXIo
tSSwYePv4fNPSoAV1DoybhlH0RWhZLEgOCI1RCcUWXJfYdZf1rzbkQZ/gIlLRngopax5/QATylup
lTCYT/RDBUgVWWiGWXQcqFcpjwXSs/TyX+GO35Gh3QMpqES7/3w21d5aPaIVwpB4G6THRhE6muvD
SaAxng9l8APUPB9gRAI8N9GDgh7mBS6UVnx7JW8KVJ81264gizYpYeHBYUoQ45AtLYsdc0DDF7OE
f8vvIjPrZxK6dRH0NX3t6xWlrzHJUZTW3W4UP/P99Ivv93izfINIcfHPp2FF399osTPLATTdKkY8
+RKKLl8GTp6krMsdb/wRQrpkLDaDTfiZMh7xTSMkuNBS8G2wqQrj2inBFakSjlLa6Xum4ep2BDdc
RimIEYtdraAtsWfclTHnOExdbmcxEp/zn8Ufa3BiE+A2YlfpiFmsXxcMmBEwZrtoFxSpxi4+9mLD
ZX0SE8TTcp+f1sCWV4/rsYSe/8bDyzBwgdNAaC9UZTWly7DYSd7kwjrX00TKCop3kl0Dm4EKUz0Q
sP4GbiscdETsmvUnvUEKBgxTp/LhThga6dVI3bZlB8EbJz3ZKfUCjhWCOLsqLH1cwkLM9YZJb+NR
mYdK3wIp3yX+VuE9y2Rc9FtI+sCiGlcS1OD4qXEUdMwO/GyQ5+ITiuEES5JpeF4ubU/nK2AyciQT
IdJs5zvIPmwtOL/kf8E6n7AJSvHJgu2UPXQ61rGRQeiDEH7OeTQe+HbRSAeKMM9sN6+r8kGPe3y2
V8Eu8ZKH7SJuavgKq43kIq1pTZ6SPrAAUOhdCS4Xr9V6T9eR9Wz0D/MBMF6hc2Q4KnPUe5e3HqlG
O1NuqhFMyPPimCwODPcWGSw8HcHcwfBVc8r+OGVLKlNjOkXwWbFm3dHrYnuWVUOapfcvfjE3OBk5
0WpEYUG2EYa2F10W0cLEWw3dBFFrOhF+Tv/WmsQg96D8mBeCCTN9R0ebmltXL6ykgPN3u5obEJfz
mJVRSc3DgLCz3hd7ORlRgNIO8g6bXnPtr3IfdynaOrOI87JUBTNzcgDqvb5yq9+91XRxg68UxPCw
5doLTszXje6LfSmga8+1kLbykA6Op7NtaZqHj3lBTEryukrWx2L4tcmRxUWFD9yUrG0B4LnVYF4D
e8D5zF/QgEQ4KfDqyEcWyGOcwzgEuX9KhBI/nODoTPhnAREdxAOVeLk/TEWXHoLVlUbDXrUBA5uu
IXf2rhDAsQ59t/qryrzD6XuqJPK7fmnuGCpCcvzPP88yhdSQsdEcD/4HPI60Ko9qjveF6Ua4ty+5
2/dnl6706TVIDRem5arw6OKT8JtPneNC8b6ChYGm7VKch7dAMpJXHmEuYRHBqokvt4hHWslA8fYP
DMAB6Jk1hEc2ZJgHODQ9SDIpdZVa014AMddsMYfmSiRhx4C9fQ1hw23WxIwNZvC4OUeJeddcC9Nx
ozVyH7pcPYOUVZamjxcOQgc/SliXD3Hmo3ljGDFGBONYw1H67GN3Yf0Zzlp6i/PTDFy+yJuDOQ2U
BfzxbgDvC873Tw2cQMh+LUH9QVWwIbYtkCqUd9yETMIh9VOnLsT3zQhSi5xF2HT2uA/kt+BDQ/1x
VOwjEWylvdGknIr90LQeJvV8qKq0TrVDwj344dZVkBG0JYL2X8fT2DN+KrHFyLKtpb78nR7VNZ+1
1Rta4l8OXQXDGFgH1H32yDRY77UUeJ4Y8UMBzC4YhmSeXdqiHyu9bww2s6XipNhgaNuPEvHVplD4
RsY4vRjB5vUPAJsWDeDHkHq9mBzaSdC0ExsLs24/0iaHYifN19zvqSIUkCP1Z0AYmyeDeVhOG1xR
+eNRVtnF+kyyKAzznlKyXo89r2z/SX5+60szszMVF5i9ufSx2QMsb30aYNJCaJ3h47Ut8Tl5wrcw
DccS/N4Lsuo374W7CgUZ2kU2AktWOyHFtDHnBtv29LDVFctJynhF/i+Al0JwTQw1jZ+vcRDcdegV
D/6/XYZhzrdn7vByL1ozk8FbDuU1DFlwUMjR00SMUzmGBgQc7qvPp2vcPEcOFzqw00d95Mlk81sP
3wTjr09Aty/nZfqJG9jPxvNi14JxgeNKYRRo07lw9ZuDlUnK3eGA6Gd580QY6/l4t0h2zMlVpm4d
JoFBA7eF5yCdHMxFxR+C8tIEc0ZjUyW/ewPwYp6G+PczORVKop8DENI77XJqPWEzBJG61T9U6x9S
o6YEFdQyk1r1bOaiEyHzdVpC0hRCm88KvVnCvuZAcnyiG9LQ4EcZjzZeyJPI4EWw0B2xJj0Wfb0K
8c8ji69h5GAkYmUqP0uqVW9FHL5+T0mrRw+xPnDCciPyRaLDUpMQ8LsQRZDgux6Ru1tOEfJ9NTYV
NKy6QntNHZivJXrUFourJnacd8adsx+r3xktNVzcEE8JxA63mfT8c4YbFEuiyacprqP0Ze84/hYI
EyMw6YHWQ2BKrw1iGg7iBarWWggM1OvIe7aNSoUGRA4dwWv5aMH7WDT4VSzp/pCzcflph5wL4ty0
Zm9rTS/c70YB373nFKxKBwIY9REZ1Zwj4RHP/LlV8vv/rsKYck+4bJbm7MI0B7GATAqYVNJ0ChSi
1683rDasvZB/nEoGf+RZyGTLOpzO99LiPKMjlJhN9BzgUyOA5lA+obMRO2VGFjOe5gKc31WabYi2
m4M8QNuBQYCG4Imdsv3dg/zvTQuX2/8mSmIUN7SrIA8/bk2g5ciqTSoiVuaHowhxTol6Bb42jvRB
4qltksfOw/QIPRqlY1nFe6+ptj1haQzpPwbjLuibbUjGUIZazyyPDZgER/UUvu9AFVTPx7ZpJsjF
hITIkHwoXXX/735w0u6jKVhmH5r0aa1va9zvHiESaMPZ6Zy8BgDmhFtDF2uJH4QOASmIq/dnnNX0
vd+jup08EWPZdGgc8wbbPFICThrRRIZwYAOX41fjqGmerU7kWUbf+PUAcahInyBKzKNt4BNscihx
fwQPnAFV4ZASM3Z5xfqaPcOJufhRmZt+6WjBQUCRj+r9dLDaDfbPVl+R+a9Y3s+jwR3l8PzTQon+
ujecAnF+IDiG4SLsvNYM9sF5tYc18KFPOHWbLURQ3B5Z+IUMbdXwu9JKFyqHxI+ib656tTw0m2Ld
UQQVSuBUi9Og12ZvfYAtl4LJtUWj7iUNhJ5pFYpPEjzSVegzKy/JpdUqDh3Brp3DEfxqu/iA+v3r
3Le2frP/yx7LUAw8XYChOO9J9veRjGpEd+joZ2lVhPI/Hr7vbjwDb1jRB+buFOnra2o7ZJEGnr5v
UUWpnQbg710xg9qyr32w1+n3V2Cv5srBtifZNMo7WPJYj/lYnoWagcF7xGbYe0Wl1udj3CE+M10E
FAc+ZpfUdPL5COEyAlRvyaY+SdedLmo8Njke4SfB/eIbZckwlN1IC5UanDOpYD30LtfUqgYA49r5
4r0FdlQf6tgBwTPklS7lbsAQqEjd0GTbePRFiiv+x+xgo82FZ4iW7TUu8nd+27F1WqKY7RcrRqTC
Yu2rF1DOPrIWKbb2Uv9dUmPmihjjnjh1QXPeyvaUWSLpS08fQqRlLcSGHIQ+8qbs01svSFNK2Pmz
QZxBTKMqRT7T28PqSDRHnooZV1gdRL634y5alprwqRlDuGbyWK7WLilO01ZTZ25YUKzPIzM+OaaH
2fD+7lzhJwffcSGDV1oSJDbl4oUjXJIAdkDssoUQ0GInZl+gox9+Jcguta9p128LDWk/0irVdQF3
iGC1Jht6S+CUUzz6ynF6PH5lcFqUQiGP4aUQi5icDFaTx60a6xhnfoEj6ISXGABElvne0Af/QL6R
NRaHN9xNecFmBFbs69Hmo4UV0y4tO+2LF4oosJnBzShvwQSQotJciCgLY0dKWjXdiq7uIZ+7CtIT
u5xh1+4KcRsHSk4GrYjDA9B4GiKr2qhi1RzbJdtoUqg7WrAppoXmiljbGIP8HPZ0C6k8usNpH0qn
VaMPNlKtqv71o/E+JZRn0c1Pb1m4LmEnwTSdr/QPyVc0GoYAGSOMn+VhPHHWf60y/5iq2Se3htwx
VbARDnqyDq+jOKtTVjL0wGdqvItpSSAHNmleYeBhWAmy5SsuQoUz2nKwm768Pw9ZTCwBBZCBn+mC
HGyKQ8kIIZjX8dqCERgj4299jkyfCDWahvwu9TWSn7tNW26BARSeuiLW7UDhC1OsojIcxjoaOJvj
E/bVjsShqtSMte2tX5kW24KOtGdd4GS8mYNrqpOUEIYZk7CWnjF86hiV8TUTf1jhRXfDGnXBJFks
UykTRRbAhn6yBbIsmf737LXe6kpixiqeJAsvli5wkS69Bf291eJsLTf4SZEHCfrP9Q/4/1MyXJrs
S95mJ/g5m+WSCvkPJybXUMyd6tCVm5igQa+aV4LZCGShSfn6cXyLm0lIdD5YYZhJ0RRw5phnZ/ur
dJeODoF/kiWcs8KA/BXW++Zp/NI5ave2/YDdUH1gMVxr+gjLohh+L1URiCigfvTGgRObhihb9AsK
TPzTq+UZJoyVrTVMQBh3YZf+y5+Dzkbbw4YnVl4a/3Z9szkeS8CoKJ3pBApxvlJV2bd4I+oOcl0W
2vhp9kqNVOhg8ZRlkbkBOehhlHXHGiZj97llFXM/Lr6jU1vOcOd3MMCPq3Tfss6zZWjEl/s1g3nP
Zf86XsRBkzW01a8P65ZUwZybSbeXMlbK3Q9ASDGMQLrkRVt0hmS2cPKhyV2wPPL6jvTOQr18+xiG
VJpVAFVY03ILd+1TNLrBk1z7p1C0KLcLkMvALtnHxAewD089XMFg7Oz31xRsIZF0wNuFnL7wDwYT
yiGTaKR6D3l58DoYyJBiWF/m4pmdVy26RPraLDtGQHHy0KcY5qHpvzExUe6nl6Pxeqt7RZqfLuLo
wvD0f3LyD93IsBVgHZO+8n4IN0VtX44ewyg2czUkex0Ww/46e3ZJSPL9RYDIabuFOWOAwIDmqGSH
fP/xgTmuCYD3EAS+cwkuOo/NQlURXHvbVtryLk0RHIBwIwhfIHO4yfifpOZAAMz6RE/70Lyl9nr9
Ny3Ca3SMBWBPxBNphTBGCsNLZSqTyAWu+S7T2irBQ5TRberg5FJi2jnAhYmDpfnBl0Y6gcA+WS8I
jLxNFr0zl+B9L7Vmq+f/xqHYg2yL5U+wndKeFeTmzjMOqbt5x5pWnwQ9CLRo2niDS8smsITVdlgf
TwKdiRzzPeYu3hyVDZGp83IJCVxcQt+0KtjHaO3coIJQua/lLr5eC9NOQ1AiZEGpk++fGEqbdTH3
GyS2n6KnECosJyHKzwYf69hT5+eZx0Uz8cn9EqEm3GyO1EmYQow3DXehI7WivmTrxxDrABxbPzoL
fivSqSkXLq9Awn8Zsc2RgcFNk6r3S1gZ/B3Va4JPAmWHE4xN58FPkhHokW1e/evbvB99ob1kSCdy
/DCFxyPB+4lM6fQVTDRl628bXChRxW4XeRrA9GTBSk4Y+x0onYZRYtFTK233ywU0yG99SGRXIES0
q6tTNjpVZ8Fr0kjzJwEcvSHuUeyXz5FBsWrDZXIQwmxo4lyQRLdiaBrP3ZnxqIEfsyCO4mqHWDr2
8gjYF0m6eUoeFxoqyWgaCDZTm6V1KAUk4uhQOaprKgA5CGkUqCC5sPeq1Fnsx1nwcIY0CTnpp662
LPynV7x13SYaw4Gvit9+k9+djUaoISCmwo4voF5pf1eM7UxMA3HOv+CjQGwKOx7jVGtX8s+b/9oF
IfXIn62WzZEzdzBxdtTGrlNw0uS5QgqUv52z9CEERGiq/w7AW/KXkR4K5J/6mKYn9aKaAS0HiFFP
l2xhfwkXpZGL4OwOm63qErg/DXHrJ2m0FW6S4ZRBKjGsYmhLVUhewvLm17RSPiKsQG+UYtVkG2G7
ciDVIhDIz5v5Q7cVhzf9zSc6Sf31lghhkCyTmIeGQ5NanWUwcwkFZPNSqiE+a6l9P55ZrguWVrZi
b/oRxlsnUjs/5KAHuNU8TSSv6xWYvIu9qYXgnH0bmw93HhmFRKmHzEqLwpGarVqNDN05l/z01UeR
ulLnnJxEw4Uuvf5eSeNpgJSRHRxCqnZ3gMcLWwosvmK8wxaHHziCdV/3v5DWfwP/EKChlAj0P8Aq
h/shmYmi5PKL/ztmwCXv+6ZntrYbBgP3OoZhXo4CofZw+b54rdlHvj4BCgMuHY/g4s55u9L4T8zr
2hrmOQRVAgIy9hA2zL0N/gqjU1BqZREfrpVoR4nw2Yi/GGdxpUuHAumLI1fYG16gagcX7+4Kp+gC
i7U4f5ScrnfJwLJg7OZOjv8W4novyGpOFq41opqiHUK4YRmWN/YmIRrhVZWFfjO5YwTFrQ8d3xd2
JocRMGd/j59X01N2STU4zg3HkrF79iR/okhkm6d/jzdUwQAy2ib30HxLXfsiNgAj4shKozKK0r1j
ji3fNXvicg8xMyYM7ul2HsJaRdstP6/5r2kwpFRiXK/JYB+rFag6C4KEySyhzISfBZmt0DRStIHN
1Emd3Vuwb8YQQNxtcQK9oJn2o0aoefJEZPX3QhVDu7cICnmebwRACa0u9iNA1Z1CdS7tLVgFj2Cb
MtWYSrwCZElKZmoJgtnR8FIanK7mlkAEv0ol8GvrqJVj1M/8eKb4c7Rwl6hOJgLrRc9XENz+qT02
JQGkDkoiFYk3qJkWLvxGDOka5khOLZRzK+FnoaCfAGNmOvxluCUbiNPj7NU24GQsOsBrKtzY7I9F
3oHpTDIVUPnPyaBruZeag4RhXWsslCPKLTClQYGbg8/pUcPZT3tZNIX2U/PiVsxy3y/ZjF9fGr9U
C68ctLzMRCzb8PSeybvg/gMp3cOWyKoqSlrjcYs/1jZLR9/LGjxwrA2mtsdWBeN3ZQsUpSwtQcv1
WQ33VuxPlW1gaVi62NQUSh0boqbAMENdSee4La5m5YL0sUBEj9VC7fB7rvfQnIS3R+I1qh0KInN+
vTnYiVcjNf4aTQpvyPFCq+jSGBX32hLVi4k0eibDbjnWlslYH+Vc6bVgMwsl1RNMb772LuVM6DNO
CAeOdAmdF8+/3RaOO9RgOqsGgJxYE2mfVo43xVD9G12kd3Bavo3/hdos4WFksjK+4ZLsaQEC6oA4
UJ99Z4zyVv1QcnwwMjRFHnjIKsWvsItwHY3C7fLTk3VAQJTPJOR/Ucc7x5qg8pbUnG0nlIgIW1Ii
Sb50Bbw+8PqwouSHIt6JPbHs0ksFn7RnXydTSukNcEJBmizjiENDssu/TPVscWJTkqfTnAgN6jdl
dchs53Dzikvvq9dVAAcfjXUhE0ptrTXKN4uQTaUVYmYs5B8bJuoglbmZuvbDzZkvR9zm+DlW8gxw
AbFrjGAOYIpEAJurxla66FG+3HhmIzSZbpsvYt/nxfWpJhN/r2LRG+2+mxyfS+GpocFjacFsMTis
ogl1P0GrQzayqc57L344ZOWX0Ow7qYralbEwvHQo9JdDiQnCQ1C22JYuwmIF3WAm8j607nK490ev
fZ1P2MrPUFURDlUxXv0ciSjlEgPk/lYPi43jtlLmk+QqkWZmo67v4C8iphgvjfqIiPuSRhh6j0qp
00p/2od5gAiWAhmRlcgzXS6eeBu9PMp0BH5Jw5FdSANfv7iX6JDzQl61A+CfVKINmpPD5taoYzOt
TZv3cVJeO+Jg7hsfxDwSq93bS0sxWXKPNnZoHOdquDUPMLEta0Odp2indDjj/XqPYFG0CfoAdEy2
guTyNCjeichwZ04K6rjG98mf4jv3K522QQ5FGIM0N1Mzzz0U9tFXghJazWP2U6jvxjhBDnCxOWKp
YUzxT6G3IV3BPTql6FoptHdX958zew7bR4Vkf6aBSxEyQS/krej2eIiBnNz789Y4HpHBdphp70Nx
Tmd2hgGkkEfa1TDFMdlsrIw5RWeRtMkcx4BRlVKYgj3ymovk3n+hFfgtEsmOSeZ+DX6qPPN3SXGb
LG9L6NQdw1ZpAP/Mb5Wu3wfhG8wUCXZsSON7dVzNoQJ3a05/Uo4qee54yh8Do0kr03KQi1Bgwpl2
9UJke9WPCQVA0vPuR4VyAtYl5MuzKhSmWnEgVxO1gIPWS5hOxDZqSoSowvqvuDs0qjR3K8P+UN9I
Uuh135hlObkwAWcSQs4so2GDptdSzK9xjFVXdFoCdlrf/Zshaw3U3ny7p59jURuF7jMH7zIwvXGP
ldUmU/fPzM4OXqQ9IoGTcnn1mo8akTAMnxr90xBJBLJ7lbg3asevWy2JCEV7k4xzq99TNtANhT9F
avQZNHnEj5Li5wWiiCE+1VSAxUv6Iq2B3ORu6oBLnxzfIUP0VqfANHrQc0APzR2sLHgObBbkkSn7
W9/R4KwW/TWOYTOUHCCtnWmMuPK+RghBbal+thA4P8e37rsvhp4xrj/T4m3NH9K9Pefs+xvNUPjD
Ia0GuKoGCCPDRQZ4Diesd0d2H9OU85I0IAZW8ZrZ1nJws/C/y6J+f2QO3BzzvOo4Hehn4RbxwFOd
kJ1qotkZqaO87jBIGSDoJdTK0uFkaMm1hPLDkNyPQVYzVaWpfKcMr5pjntAue83VJgoSB3+TNbB/
3eNfHIrROkupY2wXo6FGzVEuQ1nl165Hq6kGWsrHfaq7F9TnvO5PFw26pXC0l2UoFmlhQZx5MA5a
SqntuUleeozzTmdHr4PSvE/GiUWYCxxS0e+uDJaUmR4k1LTxMim2UMmIUpKZciaUW06S/BiJkorb
CCbxmzARD9NEQFzhZ6VnV9Jr+mttsljfWSiiRmy9VgnMd4J0GF+pIsr6d3xT3VeyZ8Maph2rrUlF
wQ3cc3NwBZsXzYJLWoRx7zMtGopCGabeHr9G9Us6i0RacEjln5IAK+Eu8faFQjaqeZB/R6dHnPFf
j1HpKPght/cNrjEfbsAvprBgMOlgYoGA1NyO7ZCZepE/MeS6fbeDkb9PAJCQJ5qlbaBpHOYTC/80
6gDs08hSBnhC0lMY7MYX3vUJ+VU5A5vbAOzqCS0HFSDFk/dUuYZolv+d6v3Y3tCSbf9iduiWNstG
qWwtVGNPHHLrVL+grFSMRR2g0CJhkOn7HujfxKlwU0IWABGRPLzYvXTlQ1i1KZSYOlsSLOHKqmj6
D2501ghgUHJ6qCj9Jq8UCnZng/Xl3UQgzKJmss2oDzFNUM4Is5v8z5KrI8t8YNMMJE0j7XGTUnKE
LsqcEElhrtv15e0v6B+za70oaqwIEWTlXcF3xDsXJWmouZrKnysXY9Zdabh4Uj8IFCgEzTK4RcGJ
9tlW23UEg1j0aA/aZ7adXsgcKlYQv6Nvii8bnKA92urzDk5rCzttJ+pVypFcRjRFJ/5IEDZJ1Pwl
yQTvFay/uSTEz29hvYPqPqTwoHYjnzHc82ITthOBPFASi3UQVn3uU6yvB+/6rj8XlBpPsLu2kzBc
ULPbzAiRFus2vGOf2VIMwF2HNswZ+rpx+mNcwBpVxx355gfjTlvFArQyDgOQH+WCKByz6jMe9i9C
0fyuHHGFSuMplejvOpJ/1pYma1zhEz/1TLGyw1WI1G//xQ7oBNrPFKtc50zyFzQRN3/YEFWuvhjF
taPy2ikMdHkqMp1t8PVpt7MbfVv2gYbudtpBUpkGxYGI7P7q1copS4+dNBspqFgaEUZNm7OU4LLP
3EWqTpk7G1BiyIOX9FEciCsr3TicTw4VfGMvUN6PUZY3pg4d9kZ8td2T6f4Yj1+JoZx35FdqkJdd
K7rA9V+fCVcKHlPK+Ey2k9yoC/06N2Mnzpb0wedn4Ujm7Grr4nisAIA2Gf3joWpbwUEvANTj0V3y
HP8Azh/YSUKNIjV9OBCshIK27/kgrHStHnSjeZRQWkbvtmohizbcRHPO88N29csHOkEqZjwd0i0W
6KvM+DNqUi+s8lr3WCP08NgDW45luNI/j7GvAo6u+Z6gSKoNLBpr0y6V6ELfQH6urpvN2tl61f3e
0gNd8xul3F/eeoPUUEX81M+dlyrFSn29hD5UEM4WT8Wp87k7uhCZUvRVJiA61j3A/E+zlhr/SB3E
5pnpEcmh6el42MpDwK80pce14ZD7fRwr/mjLd8FlzNdpCa1CQLpeEGTZsepDKQLAwdSL8PI5aiaj
gk/w4QudlUm3CXwI/uPUrkvouHUw6MGVJdEqtEIMQI9mlZKYELUu74vqzx0KZsWEqp1JWrhPao6l
gOgnzpBtmT9kSxAFOq+LhFgATF5AR2OiWSQv7r+HZUKdq2oAfmiKJ2pSNsd4jeP/EFO83AzXn2Vy
KQLlJZefE355ESEDPYsIPnb26IohSYkjw15nCPO9H5umtT3r9LIBA6VXMkzr0i8E2YxJraQ0x6+6
3foYA0UQ2CL0kUgcDg+UP4S1iGSs9E1uUGb0rsJpiulYqln0iLjDceGpNjEKY5LpakOhJikVdixc
r0sDxJa7lUvGQOig2qiq+jOSBh4D/XsCQANPnpz2aZ1I7Eao7rd7ftruBqpRQsCwaAQaFFi/6t2w
lbfUcYAUg0BzN6eYJb7desIp4ZkHPxHYc2tQI1esVGCCCQQirAxGEjMeduTLcIwK+Uu0kqnknk0o
0quqwF6RRC+KRffwKX09v2mVuvGLKD57phRqOSIDJsfhFzTJSkd+nSgT82bKGXisSwb8Aw/oXAt6
rnO7sKAal1xoT4gRDS2vv9q1JWFei13JjUE5PmxvhmNlJifHT5w6R0TzBLxFK5qd/quWOEP7HvMj
ZJ/8DvL5TR9o/8hRmvtbLqJW4IxboQGXVsCBBbkEnQs9fY+GD53KgCwi5ke6yRsoDEu2u4hDbXFY
XJajx+sdoDE8gfHjbKTD3YH/D1dSyA1WYId9A/JFoozA6AqHogOgGLcUfAXIoLepRvbmCtkkqz/L
ArJRB0F0Qph04T75kFv4GQTtPBVekUH6ndBNV7oHXrLfLLTBVAYvblUEvP9zNmVuE+njqRTc+Rco
8PX64dCbEfr35qzyifriOrwsBsE+9zajIxaU6xeB22dC93aSYqMtzzr3Et1rUH0HImHXOOaee5Nf
kTd5IYTZj+j/a+jAXN8RfXeudNbuQe9XktordOvgI5ETPRSiF9WfjpMUOcaxNkYTes8LJp4swvlQ
0rvuXKz9XTYrfknAjVhMDRxhqg6VnNysj+AdrxyGhPthkJZbwOE2mm1NT/KYRXUJfw1JOWfhj3BY
ymqs9sK1rNqi+GsI8BOjHCb6KIg+xNyRF/bcK2ggkmc1mIjwhXI42KTR5UeiLuinz9HOamECdioV
4YCKVBCbI7ADf4wUVitXFeHpY9MsRsMwsx7dUnqLzpB6odrC5hKXCp8ndnGKtu3UR469c5JJLsdk
f10JSsOfwiw2WKC5oyRpGyZyRVMCQRBezQxv6TnBJ3MnDuHZp1edlIKDTfe0DkykYGSdhalKxKE/
zWWlt11ZWcm0n1o3D3ZCdQOqrYBNQm9j15wcB34Pg75Zug0N1PU3gX/e0NQcwxdjCQRkbzNBE1cZ
MR6UMm5+5nH5jcMEGOGGYIN95RgH6kfM34eQzOwCGj4l3Krbak2c51gaKJv25pxbppC0O5S0oVhs
OZwtOhW3LdL72AZdm08wRR4UMFUvg3bDrJLMHGBnU0Qf0jHDno4b8LIUsVox5tW0AqxtOfBCLksL
n0XV8xtt5bnf0qWQtaT4mmtQwYE/AqHCPahCw5NUBaIrz64bgUC5JPfzxkd6pxpK8eucRjiCEyVu
Fya/SkbE8sWOYjXZnYIQXzr5Uv2Ur8fiMrvq9BMy5VzfvvUSD822B+KO1UrIPUHxzgpX5J0aBXye
8oOCSNzBTOcKRkqH7KimpJYxrenDn8EK+IyvIR8WZ2c0gil7NcGbbAY/pzgHoxOi4NTuwnRg21yI
1bnHdQO0187o5Ldi9/y3tiF223UMsTtfeLE7A1nntJfOMJ96vp4lZmsKBIPyaKs+tngl9fQrviNj
exB4DRp9SGkLCOCyUmN03QQbBIY+FbUgPbNdi3SonEDXm3mLASyz8MFGO/S4K+Xu0CYDYrAQ4qiH
VWwQJyawEypQnYlcCwoXq+15Of5URGf4F9QRGwBbrZ3gP46Sd3mBB7W4BVI6zaXh85teJvjOtbkV
rhUoHDbDP95Ofybj30pAbLfFdoQgkYy5as2sqP8TIaGQM5GPdILVP2c99j3Lpx31XrgV4xpGUw4e
AC1tB6z2Zznj0mOvH5MiMZuNlJQKu9GBsYP13Lk+8hR32NBuMo+JVTWMyK7Fb8iAac2Ld4ISHn7o
S6sRYgp1uBFpNaPRJX6qAATyCuHL5vX6R4nubpUPXzv2p8KHGHIpIPxXyH8T9Ds0C4BYu6lTVnCM
OJiDUr7pW6Ohr2wiXWM3eVi8qiMjgPUk1XbppA7g7xuQSfjah11iggop3+1IMI+HPTD1jd8kkWXK
xWYup3RZnmdEIX4u6SPTbPRmWQVqgCiBS80fbzpH5mRMsmj/ZcZk1VmaHokUvOtW1MFPTGkEzVsJ
dtwUaQsX3DojSSE02VwznXo+aFEvPuv+yy6p1QkGO7Gs+Iyz02r4T/7kUSUYO1JA0pRDrJkfUWWb
KHJOzxrgvh9jzNIfhoK8BR48J9FxpH/gvnH37vNVCbqt7KOZQ8on0gPqk489z3UDTcoXeSWyQTEn
cE4GqpbdE87U7AlZVI/pB/sMK11SBBNV6njlh5X7XYswYC+IzHWiinnj+zqleiKPOo5rrkHT97hf
s/ND8AX1ZPDIRxYhqynkkmaANMFyBkmRSMrVLHoe7oO1VNHfq300wF5WseA64wq0cPH0gLEgCCAq
35AK3aaNjMPKuWkYC9COjFz/1O/w6sDPaYHn8rkyoDqPngJEhOI8sUKh623f/jUIta7Lh0gzl3TD
OpgQ1RNJIw+hYQqwIgE7nqwHcH1Fdc6SN3gYJLI/Qhd4m5QlVa39UTosN1fGLkx0cTDRAlXJM9D2
zlPZEXXuSdYwioHMLHFGcEhgZOGlzimHFbkeG15J+PYr5fhmsq1r5uNUnGpjopg0HfXXpI2B9wQg
DU0kb8/elUmKj95ryy3bXJZRcaacd43Uvr2tRp/bOl8tDCYGPTiZnHTEe9G+RzOvLGp+cBH0pJXm
7+yUYR780Vwre9UHZ178yMguc3l+442CCA55MEA7RaN6EXeTeaK8mIkreeiwXtyitLYKSvyimXmR
h8OZZcWa4R9vvcrnspPVpPgnyUquYiT57MG/jCRl4rvfKaZVaUzF93VkVUK9Bo2N7z45sRkV2aNT
zvvzgImt32AAPnMVo+HYfP3O269/fShO75GjvieacwFjqV3N6e6yUsTex9e9sJj5T70xwaozDFMQ
0HYHneEHThzH7I0grJxuiZVmpqjs++uq7eo7CDzIj8Ntx8aMH/2lqnpFt63kRPzxKFy9+ihICvw6
pl7kdS3lqas7aQk99/zsr4tIXeAvvDHGC2zRkPY9WjMwfq6NKO6/RJPVcZnjVOYn9o3vumBL4TGn
7wSHCcQwsJVqtxBl36ZjxkgRZ0guUpgnfT6k8uZCXrmUXVGnndFZz4YwAfDgSBL+N2g5djOGs3Fi
sNNxUo4Q+qhIfmpFOpIkS7c89QrSI0D35Ga8tQxZOa3m1d+lBsPDBOtRI1slRy+D8CeaTnmGTcBP
+8V4xQjdO5/W6NMHUqCfavjRCASajm1AKIePqQc9CHjJfeWUCB9WCvSTTo92b27J62QbEsEAUAQF
h5WfOYdYq6S6f5jQdIuBjrGtyPGcZSMMz/kwv1dDB82v8m1ytUSKIyoPGqUZfMN6pKPtVFQWfsbW
57Est69Jua1ZJauI+/ZRCk4Q8qSPvb48uOBZuSah7yW915PiJ5sl2zHo2qUZNu7AABXVT0v5MaNZ
tmesBQepD8P+ssflyC1ayQjjpsJU2jQwoPYEq/ZVOFSC1qcz3jYU6jA+nscdltVf3u1a0jnNbh5U
1tVGzSTxjMZLg13WFX2KNCpXZbm5zZ5xEkcKZe4o+lAtY6lDYiuM8+k/M6VMlWr/8MXrK7OE53mr
J9acy/HVUgC78CeFpC1noxk2aKK3itspYpW5og3mjYMw2xz3S+UzoM/QG4PeCRgL99TchfN9XRnY
sMI36Sc9LD5uHVIdqtOsPg5k84VBjzQsCdfbNMkBF0onzHUrT1j0bWlUpuf/jzXuP0jZl+XzmMQX
VRLM6/yKjWraqbhduvH8AWR0cr6Mb6MWXl/50wOc2J6GF52MjXGzVCVFZfySy16PEAyanzmZQTXS
2jzhyB7Wud5t1crlVioL+aQ+7bXpEMnBUBXsja0T/ortvtVeqb1AMnqnm0Wf0zPwvMLlAU2HXyRd
V9e9aTaQTqoyQqt5CCwKBW2V08MVYZrBXBgr6w3JKvScga2GoP8tSgUz+ei9S/joEtC+ImHwK6lo
n67BJnJHOXhJiRYEKioYFPDo3yCPGBpvw/tAr1oKB7ahScbpDNyHV0ZSxOUPwN6PHgpgyZ6AeG+6
Qjm2bqPdW8NE5neYKc0lKvEIjm+irLNF1F3cmHy0CXBQnIw/D3AowKYo8RtoiRyAlkhxHpGqMl76
moXbRk+oAmhydc2LjtmYsMP6XgGlMUMtwHVqmQLgIsx7DqqncWJ02mmKWiseuCt3P/Nmbs3Vj44Y
9D5m9EKrIa1ZlCarOaFwlEvrF4KAMIcA60y7G447Krs2HR9VrlSr13NGeJWxVfWnvOpV4OZ6V5YW
tJNUKnyxzBOV7EEGecxwjKgPXJsXVOOnUzntIA/zKMyUD30V9yT4y/T743PvlN0PNmN9fs1Bs++K
xdxWIVvLkrXJ5R5J6V+OnjpJFUKRHQ3X2ik8HUfa0tfb6WWGEhy+y8bTVs2USG503aao5mM/gkzD
JPAUOsKswVv+2vsFF3psLm0YXXWww/nbP4b16vsWCAYiwVTGi7Qz6oG7V7Slb1s5RfsbI7MWQVT+
kRTlyVT0vm9exWxf6Zxn53WD6hPkNDN50eCHDw4OLjX7MV96cOCUP+PQU8b5JOTafvbMbmA8Bchg
hzUYm8uNylIRw38lJ0zs7FN+31pkqz8QylvRW1HywZoMnlOuyB9UVv71/qPAdVKUkOpgUF3FvEoo
kkb09yZREmkOo6dzVQEw6VMpI00e/YoxW43vMiFSYJn8kGy6CAW/JLv0r33Tih6NVJ3R7hhJ3NkJ
Khxd31NYisDAwcbGi0ovgxW6UW0vsUw0se1k07lPa/J7VXItM//oyiB1gf+uvO5Z6yZiW4xM5DVZ
yEpSw0uX77DY5YbAD7T23CfCuEFZlAsiSynoDH9YnQjyq2vIS5RL+BJztnxlstFDqbK7ZKxpTio9
duTLvkgM4OwETD2WaX2UjNcvkyoePA/x3c7nlxn9dj7gQ3EdUGX/z04nDYeSNg/g8NlWeiI/mPg/
rtOeK5ZmNHaOIDQ3WBsDfBuZ290prll0vKENt5Kp+WMo7a5s2KuJVh77c3OrLi3wUVch8Vc7TvRu
DuQ2rsFQvUqKWn+l78IZ8ln+DLnSxpo5KnYK8UcTNzdbORA9yJNLSmol1lHIw+CbJXB/VPrSf6St
0m7fn6BEQ4LcfQJhPHtYiApmUlmqI07vAGeu2GNRSAJa+oSmbIFJo4xNgyfNWQQpCu46NMEnjYYZ
0wvw44CF/3mYY0mSg5ka6lJajUa2XzQGbZEKV3pbXOQfnNwtidiI/OKgDZMYYdMGSyfNInNiMiCX
0gvYAYPOeKNuiKzweXLti2ZWEME87GMtvfXFhyktF4kTPUznCNt4RYNDpg+5REG/TvEznEcGa56k
CebX6wbLV02zIkQHHubkx09rBem079mhH4jG/uZvKI6/UD4Rm3CLZqmLI2JTE7ZTASU5DXcZvwrT
0Y9zkg6jleB4E3+5+SLm8UPQag/TDMvXyz3HHL5NBkzZfp6oYfxOT/gMZeh81PKT2J2MMixjpz9i
PtQVEOOsoJTMybTz2qJEY1raKkamK4ghKSppy99zk0JdDCmJH7jo+kRvh7l03Lhdb/Cefl9j5ihH
enttWZM3Cm7JK61yt1Tnfl4yMtly/w601fcZb+JHRI39edA40PopOr2HOOwvXjFpGmVPtGviS6Ct
07ooWR+KDK1qk2xz/kCADZffrMSRK0ZAhn1KA23ElZ1Z1U8MjhAZNjyLAiUhIiGqr6TDOmdxQK73
PYq0YYWGUpdJfPBM3myc8DaoepJIDJ8RRiqH2PXVx5QbLACXi27/LL0/mNkB+7skrRZL2H6W8uFY
ZlJpZpfHLiEPQYEC+6k25OxjlhInR/oKyKG/kiFLOKViVcXs82qp4hzMe5aCiYwe0rTi0jy6JzJs
Il7VpjRVcD6b824MWp5zz+0YpLHW6bJZctMukvY5AFgLqIuFOd7UT84tM8LaFxzZRDl5XCFN7Dqo
G0eSjme92Pbeug75MNvzcUR/Y3c/JaV5yn1UuYWJP6yoKT9Syx+MiQH5KFedHHwo7zHPilQmnB/i
P8Q/+NQJK9FQFPofw4DlNyWkl7mpqPIBYlJ8bl4zJy89gu1kUWrBgugM8IvdvXrACZf5zugbT854
EJyEEpiamfTDRcOHkiak6sSoBvngGkSf+R044L1Qk70iF3c6j5wqUU+PHPYE/yCV6pwGr8Vgy/tA
wPHV6kH+3aXRaog1GC9NRIjep0L8z8RNi8y7eV/1zXVQn3siexIz4XHTtsxAxmEL9/YqfnU/tbBC
xe0m8q1Q/0zaoc0AmBBAr6gK6yyMDWzy2qzieaBqu+vEd8RXOLnp2IxKSA7IgP2eKcHltauH3kA8
aMh8cIqF0tT1mg+eaqyfY+nuSwS7zr06M1jzB5kYjmtAMEd4rwAMDfAdS91xCA71g91AIA71uB3E
ZlkpBrScjGltuaXbTv7rfYVPMORrUQg2gD0vdE3gnMS7dbivbLeFfw4rJom3UUohHDeUWu7xV3Iv
GvdXRMc6No6dsGzE7RPoIor/UQFgYEYkojjGiwg93FVLlyQAZVmZR7erYseKE+OSBliDLZGkRlfC
q/BwA0Vy2IImp5KmU6O98X3ZoOiZ5yCyA3bBkqzOWJnt2b8pL3Cxt1QZndmlVVxhFGIHHEZkz6qO
qFdC/CW1caRXbcrDDLo7chyLu1R2vALiQ5EKqE4j85Ce1z9fFg2GhTVgQ+6ldptVG1cGJFxoImz2
DsqIeXEZjPo/zq6ncrzkv2DuGlLYLIbGf3cWHlw66VTxKHQr0KgydUuuFmvfGARbU5jx2ySOHeYu
327SbGgWLo6zDiEBCv0Po0qbWbhJDrKmNTWNboMUKC6bcfvF0ZDplYJAhbwpEX7tWunw78dCCx4E
OPoHUqHowaD72bA/n6BLbberzkme0BvdDP6AfNicSeDLODJ3wpUu7GVTUnkMGgWLdSwJwVqNLZO/
NhN1UBtDu3dvErTvlpWFBw+FQW90Eu8ui5smpwlQrVVS3RuJH8xdKaxD0eW+6Ae7wRThIRKRhp9i
HBxjI3PtHkUJtThCbTQSx/VUkaXLi7LplsJlcpFANG2qgCILuJz4Yj1fPJGFv0WV+UUzCWLy/XH6
fc9973CWonY5LC+tQ5W0oaOzDpRcPtS7rUn2A+UhoNbraM4VvuX3rmSlC6IpFutmjfSGulXdj0Rt
Lb5abi3Vtfm6vM2xyvO/xXYAMMHRJjx7ljT32jWSqV01Git/b/+gzj/KI47VkCwUFRamcY8MgX9X
s3MB3x9VQvu6fRWkEFXp8P+STFRhDwIgsuvekWYM4fuqiqoxoFGKEkzzmU3wqqrSxyl+20M4r7yx
eUw9yJDGjTuMiBxtreH+ptXJQ/88ncZ8mR4+9k0NCT3ArELbq3GOFnfZUF5HQKjGAMzkWKqvtmpM
jTUSQBLaRWhmAX9iT33IbI0v2gW3GlWrZGKNl1WVUDCBlZ3oLnCd1OmMSgEYG3MsYiAkXZM6xMIU
oLHZC33icJZEedWz/sNycFD/UYF3mRgTISlMCDEuqsbx46SJ+Ct1Hlhyig+2zmSPB3q4yW9qrSfC
QHMO0OV2q1+FKrJYuopXAEQDzQbGjUgNUeof3n2HfCuZ2HcINjpr12RAPfr1LRrRbTumym7wS6dC
lfJC95S0aIZvmv/yhUWsiPg387S8kN66wAkAvROu5ftrQkzezmF3PIgbhqLOetom/+8nnHbIyC+e
nKWqsfyjr8ELxnzvBRKCJFDZgfAcFWN4w+1aHhO+mu1upmFwNy1tkDb6y97LVlFoxpwQ+UHVqsiP
sUzCk4F2EpukXOTRWAY/ugXpab8W5PN9RD1lngTP0qXpbD7sezwp3ugG3VH4NNlbDcPLof6+xFmi
K6LOoYhSoXXz1P1VAqdonoO9GoA2skGykeKRqn6/jMSiTWU+wT+WoxPpH1m913kzBwQSGRfcRAHG
qYj5vEA9+IEEzhj8vXIqelMlYARY8eHOYkQF49V57f+6C52gWBbYwN3GRrMCwr+aDiAAmh8y5Kr4
GeJ5nUvgd2ptw6hdJW9GYdlabW6nqJtScZkILzktJIywfeqegXp6roXG16pel9JxRWVYZaUWHqSL
zlpNw2IlX0Dure1eWiQwkjvhSOjNqibJBZt9IjBTTH3S6Rk7mhVMATYS6C34gw5bDK3EfnzaWTYX
h0eStg4RJRdLrNt1t7AB+5go25yUc2RedyExHomf62gGbzxp6qUtF/Swc3rGfnnJeQZg6aZ9j0SA
SzXQCWhEomHLJhBVGOKurNggQ100mR4LYP05DGDo80F8pw12DhJBfNh4NZ3Gk1HOe/yXhJezuxKD
Tv6jOHJozq8Q7iOTZbjvkfG1Q2uchzsAtsqyim6t26ZZEH4PERbUncmXejFRfqeK7tmcN6knh/6q
ZSK223DQORbAcXNd/TvvymEZKQURBACJ6KTytWVrm+AlTiao7OOPXRXqw7CXtmrMkxpWVV47Wwz4
LBGNH6R8yj+B4BaffwqHlAiEZtxirmR86P2QIbjI273cboSohutT7/MOJ9BrLrBYkrQJTqmtcOdN
S0h3Bz710FxxkkRlDAzUnyfHV6O1O73AevxaAI5KZL6/dkgv28PempbpW3FC/NC9S1EAQXdmode8
NhoBptPyKSmUcQvEiG9p2n2szbdLi6soIqdENg45qDLGcp/k9c1Es35QnjSp2QuC3VjEKqAgCmcn
Y0v5YlDkZK+13YhQ/3GZofYocObw0ZqOnVgHstCytgpHpCMyX6r+k+1tEEwSIV8kv7ifKmNsEsm1
zt/rmOuqlQEPhL3DbLSzk7DB1os75kB58s+udb/7qUs5asxfHYvYHkq3ft73UaC2F11qA0Cyl9cE
q2m8xk/ZRSixASUNfl61XJUjXRQJ8f4m6UezHW/7Df0Bcpw0WNDMg9KcodM24TtuqM+EZ8iwuKBe
/pI6ls//+FDED62KPLRFaxw3Lc1NyV0Mg7UPlISDdfROD7n5PZMlhET0xgg9rkQ3G4bcb0hZY2m0
hVdhCqc22717nzqCDwW+lCcm8AfThf8QJ3mFa0/plmIpY21HuuZvPcYyzlnk/vvzW76CAo3YkvG7
ke7V2ZnNKeUVK5iJmR/jMKXrgnRBt8ipNKEuNgsH8xY+/BafUTztRepTOeI62fMpQYVKv0uP4Xg0
gwV9+ZFQuJrbUYn4/hMRlty+qz+hdrWVfmA33FN8FYeijYib0jRPIJvK6XnYqIJO5v6O4NQ8VXf8
WsRlKSTktQw4IR04826xCSG1GQ8oBjyR1tePRdpVJC85sJPHK4T5kr6KeenaqHGq4Lsy6yJiCZ/G
8lSW7L5UibkDGBfKDXX58UIouYsUBtaQ/x5s2HQsTwr+jsl6F9f7vASVElfF/ScXkTP2FGyGWjCb
Jyuagqj7+ScssjHpMl9nUqM34tKhBnWuNYQbeuYZITufh12xiotYBfhtltJ7ggBc8V+n5yMyQFqp
n39qNaiyu1k7yHjbPlMzsWvaKyfEWjkSiH3rk53VtnqxdyHHoYDHC9qwY/L6H2ZLZDnRd3C3gnra
R2OFG08jBfD7awhslqHGRmYLErtowbS9YraTtKPCcMdYuI0488ZIac/8piNw9j53ikYwg8N8uu4o
Vkzyj5yoJMaOcuQrZqo3qbEwxlk/3KSElNQW5fIAA228711gx8VJag6jz8rTvIqzdmiTTNFhS38c
cKTPaz/8bJpiJJf4b0v2c+pEfh1+aGik8DTSzMYXb/hmhmw0DMgv0FlKQVIpJon6UzTF3ITjX75b
3u7f+ajDUQ7xEuxbPdLqCSi/O0gnu7ZLO/19hURR12k49xQ3wwURyYEdw7HczHi7Y2SL6F8X/XHA
QycCB3usxsne96LOx2qZ/Cen6gb5shfFR8UBaSxay94oB3NcSZ8GOOWqsI6QEd/ANhFgdGUSRf+d
HHkH4Uz2ObJf7KAlmNrhsI7YiZ2aYyI3xdlu1oFpxIHwHxSjU65Xk2Iih09a2dil+LBG7UE6CKk+
AqBHx0+2GyFUmK13lg2Cu6IQ2Z8gTW9v2OcmFS0P4PgOI6bD0FDTb//clW3+qc4NQuAL/nVYOPlw
orlMbo5t3r5ofilr4MbAXuaSiWlhOILiXhDmQqCMfdEFKc+wp6EbW63c1QeBe3tRLx7xBIglSASa
5hP7zfaRNz4GDV7X5x/EAdk5sa7Ll6Siw+TE/jaiTV8s29HAYUD2sSZHDcTS1knEkbA4Tdn9wwTu
DQ4RxEy+3+DcMO1Yct9JPKOcZNnkY5kVcjItneVtB5p8qymOpAHvydtldSPGF0Y6CJAYxMJLA/2V
H1p5FwFWLtP8Y4ecrddM0ZAbP7OL43yydQMDGINlX6vFcFMgsrYLG/Bkf35Uj+su/rJ8QKTcEuIx
aWkzyja46qbEF6fqPp/D2v+jHN9jJSUjZ60U0ZY+w4lDy1VqRSh0qdxbA0ils1forHfHknwx4o1N
LGOiSlxpytnHD9LZ3J+5gWutUfz+is3hLxoaT7v2NHKVXfz+UV3kyXt6j39NBuQc0rq/HsKGExKg
ElV3W11FR6swnn/wZ73m9bDDmCdoWuSc0ffOqvLRQat++OEmmciKKuvt77Cskv9DWOIt61DCFwTp
WO0RaOrkGgtzhAGd9LIlAO8q960h7PD4aePlUk3Zdzo7/bvvm6cEqFREWjfibWCRPDOjFCyJvx/3
rH6AuqWWkHa6pvE8d6BTAPOQUoIkIpxGN/hYwQIr4aTQxexJnUFDrwrOHWDnP+cQ9evhZeNxy4vN
ak4h/7LHdnBSlnDGkPSRHBvqzq9X2gbtM6wFh+U2FLx85IVCBjPlorTwa77dr35rLSb+BNxwpvpc
r7KTV/k3EoitWnBz/noD3E6yCWE5NjyNZBLPB2qe/+yOjaf6STvBjUL9KNYLEVBWnIr9WUogDaom
G7z0riQNUO4vlkAEkxFQfgXKFe4j4quxfMe2Vu18YIvvH2YaffVp4AYPGYF73xb4qPjyjwaJe9tf
BEPOSh5tOhscd765TAM73+ykGQ6QgVW2VJqGLW1QD3slQ7LtLpePfvnvEsvuMaw35XS1J5SQJG4n
QD7Y84rvTa2d8QIC6ITcsuU6trHtU127999En/jm45O9rj0oJb4G6VlrA+uX42p+1i+wIy/mEmfA
Xd2DgcAPH9OA8CbrkxTeYYAF538er1s9xM4TBLHSS+IZXqroYTdxKR3vDqO/R0qUXsI9ULzmIt0h
QuQmpP5yYibmo1ODg2KvhtwW7tnVIJ3Wqks23R9IXf/mSkmT7RWdzVThKSfpyGIkCIj0yXi2osye
VjrB8iOvlXX2DSGbE0tntb35LeVregby2+CNULdIU8+jyBRg3w/Pg5boegDGCkcetSvpcPIHo+nh
48oiUwEU6qC7zF7yQ/PTTePNQ8OQTm0EtHSa6uA6DJ1vEHSkEblPtYoixcluHlJw2oSuEW+kwi3Y
N/Q3wNcdy/ipabe3P8tJ9EG3cP3bjNWqpsbOtE2qykNVo69Sda+UM8PJPrmnGrl2TNbfBMyMEi2B
e7h++YDohtOdj3b8UqlYxLMly1k3imyUHsytNi9A2c5Dw2Z3CAjHdLA0dRrNHynBbiVDF28WG3yW
H/aZxZHfIt22qqWcQeVzQg3951jkPbRbUWsJEEtLtSJw9UmAi93Li697lHs4mbY0hDKNyMtmmD60
SnL4C8QuxwD7J6k+azgt1U9AJXH2GPyMykOiMwWfHU9EazHZ56k67hUpLQ+TTfymqUMi7F3CDgDc
TqkEWzAMEkx/GdHyaYx3RAPxYmOcRkehn5fPrAON0Lw9MQPta6DzXgk/RB4giNuwBiqm7LNCAnUp
E6YX7Fuhke0RRoab4ljpCxitLx6JEIe7sQmw6O1V2TXcV9rFcLG2y4BVbdtG+HPsRbs+9Ez/JJb6
l6U7MfQfYzv0SJLv9elUjl7RJFmvWpTzxQtM1FQzKzcH2QbhZwijZLZvs6bezyMVuPS0jUvPoGq4
eHRbWirULUNdmEF6duCUOQOIvQK4nlo2hIUL9JATJzVz9pwKA1OVENH59tjaAYqH0LnfLTLRcZpx
DlF6Ncd19szJ5IV1L8MR8BUzS88xgk2y1IJ45U4NZbcvYa37+feFNVkOEg4c0FMNrB1D6VnZk7TY
lSEeG4mZv9UbI5PZiHWdZkgMZwp4OpSCXu/MCo45guMfohXb437QFBw6LoBHtZkH3KLFN5tBHl4/
sBqdruWmR9gkTDDzIcgqZ2I2psnoZIl97B9Lg8PO4SyFhT6d4c9R/NeMkmYa/pDqsC2E5hxoTKPl
zWD34QzpiI1sYkaSvpNH1oXyTKO+6p0Nfv4FTiQxgwhTnYUeOh/LETdR1n0ZsjjaRnBlrSaOmsnF
BpFOzQix0uJJSsHBn87qp8kaVlq60d5snOwDFgS/rI6GYQQS/T0o4j7qPHz/WSpDsa4vrH+H0oWr
no0J/iJDfcHT7X5RI7nVlYvvERLoUvuGjPVVjrbKVp0922C/O5dGqWfB342FRIi43+2m6iOK1A7d
cIPEKgk9u6dTNo5YdNL/lXL6SeRRhG4EY1WJY1nQfTShr3D62G+sNxOSGXfy6E93gdhlAT1hr0qM
4ay3vNDnMrCzV/pwyETnItOSu9QKnGLyzNRFM7C/2se1Pb+elbD5P3I8yBnn1nknfG4Ycs2xkwZu
JudCtmN/ZD9k3LWvXnxaDjs8jen7I7q+EaXMo++w249jYXJkTdm+Vb+v5S2Cnq963tqwLd1wK3YA
XHIiFmkoUpKhxmGXfJPZSWWBwweED45NSbfvRBcQI4wGBo+TxCElgkOUrviG0KQD6FdkRA2DIb21
W/6vHvPL9S5qU2MhXBAgRe9YcTBQcSSrgJaU/mwBef4vHP6V11WBX8Jd53Evy0SatjNqr4YJ5Ysg
R4HyxHsw+ZQ3BzqsusqL6aTlYJ/ff/q8TPLxb0G6ZjMERetVn4aYoD6XVTtCASz+PwTJxA7e7XjO
bcoxfNgH506UJR4n0Ef4Nqo0eB9GF0Rgt13LaE3ysW6VEWCiCgxQkhu8ZkkR2AEfHBWRHwQcEB8H
nk7DudnOjUKgZafILUa52eQq3UtKMjYVWlRlkjQuzzniHyaWrdqaO6cOj3BBcnnue58yVikcnkSd
bIQPRPEbsBRSkvVqYniUFLAG2kuQptNeC8rwqb3lWfyJ+iRx74d7QtJbBCI+cK/qkiiWoYwdfEqw
vM9cLVNXCv4op+KwYiC45JbG+S2cjnrnVC17hJpfBBFM2TJAD2MWRH9geY7BUbkg9EJ5q54USlLy
IJK49RzLPuA5oO0apFDyfvQgqi2r2xCQ4wG2IyqZu2Ds6R+EwuZoBVQKWjgzMbLvxY5CmbK/xw15
hwFcvmGZMyrBYotHrHw8isDbSks3eT3ntWNzDYgY0Ar6HmsI15ALuGlrJAbFkUGPn/nvWTrzYIYb
8BGrvzeTGKh2TSHkw11Dy0xhjnW0YDiBCG3iTydBw8w3Nuqvc27YxsbmT87MH9TNFZ2sRTq2SsYz
kpP1y9ZoxNrb1JZBcK/jxsvsL1ZsiCX2zxKIypci2+WNkZEE3QP5cDofYKXcB8y2v25crccZ9MzZ
F0q9w1ALC18OPrcvH7RH7rXWTkuTrmS90NbR8nUiG2B/EjyUDw50S6rZ6P5OAZUmAKqqe8oyttWC
gv5wwd5RV1+VaMKjSMO8q1hl2s8SiO8mHwy9r+jT0kfDtSwqalBmwnRj0f4cWPnJJiyGHrzpSzSo
FzPwumpCK6GV614uiZYOUoGn1d2k5p4wobgDu7WEFx9bKcWy49DNqmZZK78DPJYbLdnmTN/+4twQ
GnmQ1gAn9GiU/XJsQq0W2YDy4jYYL+BUAaioQ6fl4/Kn3KLHo2DB9E2EwVYXHBoS9HOQjJCtUHET
utvCGBPnMuzih5CpyhTHZCuBQLMd4y0GZttK+eandMaw+MGtG1mZhXRKxzVwiISTFT3bCWteQSgq
c0j67gg/lcGFo1VytBkFpJVpbA7QXHiI9JsmITqvXOC35A3XLwcvySgYdHVU4bWfqjp5CyI5Qb4i
ChTSe7A3tXakFXJEmQIYTQ1qkSouWlqITGdNcg/unTy+t0vRyK+Pay1SNXWgcCUnuy3Ko5g+d7mX
arYdvChpTAt15OHxOg3OlFT/0ii9FZBIShnd6oJVtKsFQiQwWvmRh1tnB8nd1KZ/ow/l3tnRJn5f
2k0DiKmAAUmTLtA4MgA0zgDHxS/bAdxveQ/Tt4DVrfA0w5wJQzThRO6vmboDvbgTUcaMmAN6LclJ
HhqcIokAYy3o2l/hpBaFUHjpRBpwBbZp+ltQw11M0ks/PqiLbIWPWT+sju0NP7X42zddTw+ZXo1f
nONtcbYl2ev8JxmvobVtcuVxnjcbAt/7UC8qm3oKEKzppfbN06YhC5a9utXBg5zXyc2SIH5ECJgb
wFs750MY3p9CNFPuWC42pyszFuEBJSRTvbPx4u3wEbEUaTVk9jWFOI4KcXv5kYAYwA1y40ncYJU5
6HeX9M9bBti3ZbI7L7PzA/HdevZOQKH/xdigEszYihiHOc45sG+9cC6TA5v0WIk4imvciNFP3S7X
ghFe2tOwNHhjS4v1rQFnkGjbwXpeuyplV5PCgHRtHjS7tzD0TMBrFHHlrvSVBhxnEHwSRu+K1pmf
L5QJ+jHv1aeWftITBGyWO1pUVVcaYOhNP9m+6Vav7Hb4TZ76bj5sA2xKDYdFegjoUyHY45xMBRYo
MeZ9fW8YyHp8PFQjPwOZDM1cSmcJdPgRBXRmGLbqVV1I1/CdAtQDW4QcGZtw5pbxIXAnDxxKocpt
i6LIk0XuPrj1L5poPvDSeCB9NOpIUxfkUXfPxXVo785P+GTTzR3sxGfsEKXbbRREkSm5ZIOYus1k
m1FUk1SHKNXECobGqMy4871GRN4royjlqJLplNbcGkuyubzdhVgxRSioPurvI4IgqY7Zjs4pj8j4
rbf3lPvvgC+QQcNGk59F/VC2gYx1faA45IeqJJKr9fogXo4fIRgAOeefnysWwNzhaOOjUeSBLXvf
gFx8TMx2a9yuqwPNn8c1y27UEkEbEU5Wz6DFyVNnC5l1A6eN6N+BvqkvirKuNSAWKddA3QF/0JO4
TNfz0dYWPpbap4cY+0jRb/u6Vm71zk7VN3/Rh/ZxvrYP6E/IE8imVndHOdQ0ZOP6MChJw4Gkq3vb
OgZ5itw7I3St0aawAJwg5o1ryhPEBAvOWRWx6dMtqRRBurUi7LeFrc0T9SDVnBiZ/bGOiRu+xvHB
/6BUkL0FNTWYERyyC4rd+F8CwKY6SA2eLr26SUSo4M0nb9IXDp5sK8RsNwKd17zOATXS2TorEaME
EQiMi5QWj3QBNQEFdoyFBoiPQw3Z9MeibfyXUq2ElqgwXJd+lLb2PRIYtlXm9uyAZxpy/4WG9uFN
Z4YDJJCwW5CMZZffmSJF5E+4yEa1DpGTjRhdu5LafLhVw5PYpcwyqoDbU2WCHtAVLeqNkK8kIBj/
0wjlTf/n3L66MrNCWrHpPEUGRFbfbEFjwTsxDCVczlYy58iWQVOriTlXKQlUdNbApV3VXztYyxMr
CRydUQsr1/Iy/EBN/Hm38LzD9xK2IMW6KpFBIx8UXsK/k26xbUxyVfesHQzdS4XxmKWbuEEjf2CR
GxaEBqknImMKhUIpO+MDJaahtMkHe5d1+f+mZN0tEeAvDqRJk/wM7UtEdkwESefJdnUAHJ6FnCOE
U9Ef77buvIGVk38QwXaJIDxFqKbTnoMNl4lxEvqGQjFoXIZAgAIGt9zdKeAnjoBN8Qg+lyZUQk2o
ykPoz/TtHgibShJpY2WwRV5SS52fgJgbhuevvyZIhYT4MMO6G/AK1CeaYxqP0OIJo3f+6vSrCCm6
5t5BZhSSmaUSO3NM2+pHRvCBK1J/1YSR4npYRsI0q0KbElgGRiNBCrnygWjqxhA8tssqJpRbSHW6
QXkm5P7L6xEPQQQ85l+IoXm2D3iCLbUG5WRzdt5iJtjo5zsHdWjnb+btSjt3OL8w0mIqhcSgqd9D
WaYsDieLby5DDEcm6hbT0+AdeNBQ9yA8mTE5gPTU056+eoZAIhy3pGi4iA8RrhbhXjEhx4kQwT72
zxo3sxCt9mZAvpPvPRUYG+DeldG01K/IXUoMVqbsJk52Wsen3OlDdW8PsytxDQJqMwrWz8KJgPvy
O6mW5Rx7mjSiOvunesUCH04aal4H4rCQ8cCIcKmYTIXMrphJilMRi5wpTkcVyvg88Gkyuozf3xY7
spJE8JBIDryhookqGsKbBxuOc524PVNzUeF9Q2kt3POLygtToeMWpiWOS5Ks9avyZDgT/OxXsYaq
Oy0ry3Ot+/XiAxZmNwN9wZFhMsLy2NJqNHXpCUdyv4mlATjFL5Gsb6c588VweeHaJu1nubqe/77R
5m4KKZk/HSbtAMk7u4/VqpWpnOAJof+zAY/mT1JfJksT+pTY4mQ7R3CKzn/z68gf17qcK7JTBkbm
b0jvLQTHYzDbclNHn2wqQ9NWbuWjpzYuEiPhi0ZYp7EQc0l6LR/SRUoSKlP66heHcJttZOXoNUeQ
TCFkTZ34yVf1wCQIHQYEc90fxxor+yLF3IjsGUE3/ISO6SaXKjHgDLYtHoTgnew4Dmv36j/m4cys
+MAUgj9LRyXsl4Rwf6ysHlPrKfJrvzUogoB/t4fx56UjuPwxWOVkkPPmfkqI+iJMPlyfZOoP0I95
qKlqJgd0cSRjuCV/A2zrdKUCnOu7IDdEeX8Nw0/e3n6v9AMFBSDzZVnMWim7PqVtLRNOM1MGJSjm
6pTyyGDWwJw0YRjm1DHrc/oElwH4OyFvxHH5tqCaTMFVK+aT30+y5LkDWB3xKiiLLZOZD7WOF/Iz
R13W0x+p9V3dTOsjBHlhyI3zvqRi2Wil/f0CXIdXvYCh1NTMzlnlE3RbNWxdEYFLP908x7vhR9KJ
lbGs+wKVyqKtpZaaPSIPDDyfrCslN2jn8M7HnpDhNCNRts9CQ+PBQL1eODFowdupopZu8YkiQTE9
brTSZscd6JHk9qKjuUuuU/O5vBHWd4hwfFGpuMc7V/kGQN38pBMo3CbIl0QWAwUz36yv97JySDD6
/5cdNCUfyO0C/mD6lAKlEiyqLb/PZ93hzkuk4faIf2QrrGAQ/r3Aso7CIC4tm+woEQOWO5fauc3H
O1xG8f+pr8MpA72uiW4h++cREgVctfmzJfHLmdZbjtVNXMTReeKWw7kGjkyJ8Tr/QOnxtZpOSOC9
9h9Vm8yXdNybu8EmgqSgfkquwxMxbsZ8xwzGoI11rAlG85csU9zbUVijRGGW75FSKOBtbWPoFpND
bbaNvf4MabGRZcYDCqLSM/Qk9eNPYpWPbgcxfpIiXsiQ+LLOQ3awromrB4QWThFV9Tfd3tfL/QQx
xr7T9VLH/rFb0AL2CAbK4E+JNXmWPZCzlMxFet8IlfWH8ndmCjjxDGrPv29MxJgrULi3awPfcqqX
c8cO2yCj2IXkEzWJcBylCYL6BtaVRz/iE1e1uxWM3qs0K29Rq91mG6ORCBqfMUCJPEgoTP41KTqJ
4t5S8K87naBnKAHJ/Bn5jbs2LqcVg2tpmz1bwqQfy3QIXZP3B6aeLVfbwmeDaZBJLmSQHHuK6ZTc
Y/f3phXP1G/cS/5dKKct25hWaKTujgYASNSd3E3vHYoNTES4jAh0e31F9zoLf6Bcxx/CG44wZbss
5h/tKGzhgk4LhpFzEpQGwN60hDlqiSbYnX5S14WoDd7+7e6WX47J4faz5WWD28nUh7Wf2omwJWkR
PKWJmgMzBwopc/lrkY6Lj8DP4hgS2qBDx01dde9Q1vz6AntNKiNTdumHeOjrb9sNpWGXzqyNap48
SaeJPi7uPOqe+AubV698uAZzMpoUyl7CnII2Q48hnIg2AxB1c91WZ9qvpWsSoF8MifZRpt8yZqKK
uxbAh0WMwz5BLF82if8KA051nE4VEAQKfcslyAwgh+n4Q3ir6PrLKb5CYKMysmRI8jEbpRRq8PKL
HTfR8pN+w2JkvnP0LaaeRfvzmK8aVCiUabb1gKHbAENBxzVzh8OZwQEHVkntP2cz44hxyY6XJ9WK
JAxQMnIjO75SvEOr4Cq7eT4Mx4CEI18bhbP5OUXbYu5t6ZU6g4883JpxlarB+P+mPovN6uQXjzDT
Vs09eg6wtowdm7FhtTPHRLbB4Xu0u4pu+0TzY6AVv6zOFOmj1BWEBlzJtoFXsNqwKE4cGFMfO9o8
KAOYAVk+jsnyVCkgjj6gEjrHNqayG9hONv3i3gk4+cLGVW4RPozjkcAcmewAeRCqjXm4iNSGKBqV
/Bpo65l3WhL9Ej/Ldhve2TJCsknwbmO9/xXLw9nvQ2hRlqPIK44diCdnb75U7V/BgAeYMkXfF3Bf
PeCDUnl6vWRpJoPA2r4jSXDIny/nTempEboS5pm8RXBVlbE/EHiYUJR35eGk/03QFxYsyvBBEg7M
DxW1wTuiUZAwwPc1w9qa8QwwiPq5rNqU30E4/4BfF8frUdm29P/n1ZE9LCr3aVpcKE1G63cGd7uG
X7hBQ4MaleD/H70ofe9rqRl6AVkPsnLXfNuD+dUCQ3ghCsdxICizkMsXZ6nQyQDsr+5rfHto9GDj
nskN8knYokEk43vcJwZEadaHnVqKhAGXx4oEfKcWAwAvGzTSpADpFgFl0eO5G9XBSnnA4VEuI0ml
pUqaOnA9NYv5txpC1YdNsvSwCV0CblGA+AgbPJAWETC64SroDZD+iilNrxBwsjPhQCxjml/a3GPA
nzduYUCH4QXNWxVB+e3cjcMvCkR6GH3b0YhJc7cahlHZNeqem5UfDClrb00lCXhMHjNrJBFsMhqm
EU//tOR1OLrQINyq4pN91cP9iXQisfQabsFWh0PLweMeUthtCYI5G7Srd99dqiNeA1hWhOakhAj9
KX36HyuoM35f9N5UQIun0JBz7yq5JDzBNjOTbnTw0iv6OuiHAQYllxMaw/iQm6YxPOvFGr/C22Fl
yzTuXyHLcWnWUTi/C77Nc5J5iX/TE4M+du1HaZElkl2LNT0Iqbm/qjdBuVgGqRuC/CV96vq0gbPy
aDPYqNUKWJ6fCUdTnaUquoINb5J76GV+BTORWu/JUAWYV6vbcA/ESj4BAF15cJbTqnl21ldurGgR
1Pf546uihWfUq/s6ITo7eMD4kf7jq6rlUcNH+DGKiXfPQU6LHMeVdoOLK2bOOm7E9dLfAofszmru
h5lLNZO8xdZarnL3c+4oOHHCjQrwjDTl3+hbDDk+RzXkIyRb+FAPXzku0+px8TdDsm+CvCsM6I82
ABviJSrkwN/D2Hh26XyDcnco5pMw2EmJKvLBzZEJ90BjB99oot1B1PrSu7gEYomsdyJX34IPCAfe
pmin4g3PY/1yaFeogaHkPgH1b9Ib6hbuAF0gZNE+ektEKlsclLulQ7732Q/mUf1Yq/80AiQrL9xZ
lEmwkg5Vn+ybMPWr7WH/MOn+SSgeF2QuTgIwXLQSSMzqPZDGZ73hwZOK+ruWtBFR/yLOFqVzjx7K
fTtg34eb6wyeO94MLwrqy6HxLNs0k4n2mRDxX0CTLWXVjHRHJonqEGeXZi7hVTFF46Vo2zXhPwHC
8D4A/WdB0JyWYBevoYaaWO2tUSHsP2PPp6ORGMRpMBn5JZTCRnm3kP3AWUnb3OiyI28Q135nSgx2
jI8eiDGfjY5N2/8fE3VAE43qKv4FJtv1/sDRiFtQr6/Vx7UJprvdy9HsGwB/KRwUdhCKFREIsIwS
GG1pEAVvbTogXQnADkTOb99SNfu3c/IyiQrqraNV8qNOEFL8cxXBfV+saYWKxPS8aZuYV6v1F6VX
K0y6OlhHdst9HF6lNS1EhMILMDxbFjbJryv2NTo8C0+yt9tL2JpUlS58XtBGvom0bCJ1quAWtG5l
rAslI5TnkbMZ6H6nAOe88iGxEf78eqfkDKCxD8KVlhw59jcRnX4OIhIg0jx+ka2Sg61ktmLCRkQP
9Lz2OwDPwdvetmtY0xLNQZk2YX9xMueur/d1bsWReW+RLfR4RxQR4DtnOUak8QFnpdP/b2h/FL85
ez+PrH46+5vUym1FfA+FnVw4teb1GV6Y1zVl7R5WhK+/KNL3eKSDKWyjCEdXUZlHF95Z1RkRYJIy
Mj4qWTmHZJhwxJw6XZXfooyYE2L4c+YJW7nx3jhva6i5kfl1fDbCDODhJFrXCQnVi3NYKODm74Ox
aESz7XLbZ6E/HysSg0Ki1aJOZmeztVE7d4FW9rho8Zby8lgGewaw72IzopYWV1ktmg0RDK55Sg2q
dnylpAGZX1P0OSFb/y7Q/GKdZbZwf8WetELtFrQeDHYlvm3A2kD/NJDEKI+ibl/tdqqCr/cP/Dny
VemMumfO0UEO8W3F6nHubgzseaDvt3LgH9bc2uGjkY5coR705jbHvQZbFR18rXcEr1Nv+qbNZ05S
Hqc0pUjzgG+r/vkwqx+RBDr3tlosJQY7KaCyN4Q5jFeJPEluqXZ3UR3tezt3PdJ1nMBg6+ikt3F5
VOwoKSmW+lkBpG54YzFW6Xr3ALXdEUNdLoUzOilZFaFlhIc65M/tfN8ItByNpmNwWalVohJKKa3G
WP9rzw36zJkjrHtOzLBduWdiz184Pgy2r6m7PJyB4+5vsKj7hTXCezoFwcNAirBQ3XIz+SXmEF55
Y3jtCMbhmBzyTI0JzwhuDF+1xBBkKc5dRkYw8pwzzHqLgO9w8cphcE//hBxujPjpWSlgkz0WB2/P
jdSW3gUl5NGvMGLbkNi8lKwecBtTiCzHRrmsFiF77fVRVLquBn2ty0CPaTFVRbJ3/q+KJXHGUlcE
BLESGoJxEhg1Q6nT8qFImP4TZED0PHuEpT17CpJ6PRJS5ghm2pEu7JD9N5xx2/TnCJ+9C1LcNqDq
xB0aAGxvKinGRI/cJ2h7WqNIXXkCqBlkG8IVxK0opkdj1aQdPa50nnYF6xGIwi0s2UIb7lOsAVrr
ESOYHXYEXUNJQqrzJS+YfobAlphwZVmh8bo2Ww/ylr8yZinmZs0eKoZ3ZEx699bqHdEsD+/mJroV
BiOUlGoniQPnpuhxD9kO60Fq/ijnHPtdA+cHQE1wWBUyF75Hbi22YJwPHsan3oT58SF9nHnlJi6W
m7R5WwBerxCOB9NXloV/QUlYjELfAfkGZWuJEeSv+HjffR/nShaW1CeRYpnoRt6DrNQkcJQP0Wem
4Xnz5AwMKxXOZ9ld9t+PFmi7AY3B+MtRg5Vh/7EmxD2YeGst8/lUtfWhG2wiaUwFX/3MI4xZwVcn
xOwgkPw8M5kRH9vBzn2vG9tGT0/qCPH4hm90Ki6oQkdvRaI3U7DpDtviZBSQ9jzIB1Rm+MCTaz9u
mgO03yoBxj4cfrQ4ZowhCirr4aLHxyQvanvKuEXM1mpwZajrLE1MdNFOsmguNgrgXPpl0jRs+cwc
5s+xhsmzGt/5JcYBFvZANRMluL/PYdsFdqDEmwwmRVWGI9ki3WBLN2NmoIw222Mn3Jvx8r/6LkkD
Nt1TdZKH7PaL/ayrBity2jkLiImKE1FX/uDRmxk/UXC3A8tdbVxdoDEzTQPNVK1k1l4VVbrX5Ekv
TgScZ2mjm1i2JA9tgwlpPnXD81aDil27x2CHnPK7wDvfTKr0C7xvHkYd8N7qzYeXK7+NBP5SiHYo
SJOGV/zjW526sSF8s5nUciDWzxImuA3YQUF68ALEZpCAxl8xUXyrgnSFoTBSaRLm+k4ujYE2wW7Z
yDWm/62LXBOpYZ7Xy8tjMFccUlZeKA3gc0dLZM71aGZc1XKdY10NQ4ystM6ChOBLOeN3laxx6cqp
IoSnLOuH3r17yxI0/acpBhIBydrgwEKU9qevnXFQPSLgCDWfXPNcQi5embdHqDICTZZkGOPbha7L
aIkeAzyQM8V0N56Z1RVR5xAZIAGRM33hfY3cBYiV5QVrFGl/gtcUCha3+LXIlXVMs18EIPDQEanw
vYIQtubtzZWQWXiPCwghPaBHZpBLQPRZXX3voXm42BoQ/Mco9kNf7VXGfuqePgEGmt0Ij9Z37GKp
SuYKNHEyWszobE2oyb5FucaX6gnyd8htCQDC3ngcCZUbdJ2PSmpv+imn7EG0IrybPiQboglOuPwJ
6169t4l6vSVTdKvTlwVnjoZclDlFUk/9hCSuRSlLeIgJZT4X1qyGQN12n+++9FZ0LfCYcZD6UP4B
XWX/GN50NJB4XnBr6Na8ClhW6KM0DrbUlEaItzN5X6oWTg28+y8Ans3JlvcohZ3cM6GyLKEG4cJ7
/0nO6dL9+tUdWIYMkKPZrNhtgtzYqnj0mmhQeQU3koPw2+4+aklr3IcbOQ6gupG1/Ia3gpUAwHBt
KR35qGsp5pqHQ4uPR/5Y3BxtwGd9JPS01/0KyzPsL3psluw06Ruw7AUI7rgGLCfPEtLOr/Y1B4GB
eGXKNUa8u/yGWeJ1/EK1hRbOdCiNyjEldxPY3lJ0htjXDEzVU05BUoFU+EnNrlpL/nHl9Qf3cryV
qhK+ySy6LBydo9r3P8+0WbP5+uZl6lOpwHL6JyKrTM2RGUM0BH73oE2Uwx/FQKBt7tDCzmFd40IC
PPw7XvX3GRan+/XTKzrOW1S0HiNrJwp8IvzNfwtgZH1WCd4oSh2TjkCoHhJKSXQ6J6exeKyVp9pu
ydFUk61qjhegzTqWwmX0BzjP9CaLcNgO5RLCj2+cNF44z6DWryuZBm5WKtsRNdEcvsFhzIo9kY+d
JWBVWEWxgtXLVClt63sMsCFkAg4wJlDje8po3RwUbvrDg5hVjLqFj+d74O5qI4tuXBtsRn27+BGo
DG8m6BomNC9qapsHUnWfeSPOjWXqTtZWVC+qUaptuBsocs8Zqp0+vH/klFr0YcS538HeSzgJCo0S
V9lx5ev20WwFyUBi0XkUbxxiRJZgRFX+WwaWQBDPUrpFpN/vjV+58C07K3SVxeGEyF9Fu1S1W3zY
+0h9py0oO+GvM/V7ayZg3em/udJw8xVPq75JLtM6SdpXpsJFg7tDX9Vx1LmWc3Bi5X6U66iCYsuA
2lqYu7UE5/xCgUejJLPA2nmLz7VnLYt3enezq//Ane3HHKsGh0M7a0lTN3cVp19ga656uCdt716i
3NggfM0jYKol/cEdFxETUb+ap4oPrqWIzBuHZOjq/mV57EZNwR1Yhs842+5lw/K17+B+zPcO6MUD
ZuR/TmRCLx4C8JPmwUDb80UJEixGfaapPrFz5wWIcAeJRpYKjmFK9lCUCiU06RRGKAs2Eok7BjYx
V5f0jz2YKsjBgf5GbDUiF+L9umwO/Pfzlo1uuRjoya/TABIom7PLPYCmOnPvY05GzsKzoLICqn00
uCh44rLOM255qdWBP6HPbMnUt7RP2GkK64/UuUgFW+d7tD12redCuJeKwHjNpuxTOPiPGAWt4QRu
3xuHdyHZTn3WJtgxJieFIo5yjDNbtixr4DvtjXUEjEgRdr9yMo1AydHjMpQrnSxrw4x3/saquj4B
L8Fj3/QWIWeF6hHMLbjndOt/0gkgPdR+U1xaB0ICbqAB2juPd+cVa4gz7jZ0xjRXZnBY3TDVUmy1
vDdI8JYeE8tUxxYHHf2HVAvznVLFVlDhjwBeP+No7qWiXZKlQWpHJOKV3Ucu05ABzNmchfK0boXn
whesY5ZDTDpmQh4jn7AXYHHiD3ddREKXL7of8arcdA14kX6n4kgkj1DoA6Qp3KXWwibPsp6GOMTr
HvUJ0doKFVn1BpfGxKxKDNn1n/lUsLwQcYukylrq4QGXF35G6AB+PzKxxbAlZ0XhysBPLHhcvx5Q
l9w/3so8w/g2KNTaTt3V9PaL/bWWX0GyHL0AmF3JdskClrcnqIHTXXQDzRHn5ThCF7qL2Vt/FRHC
rtYfvUdGxn1EbVro5kSSQk2mqfnk/9CmNqasVNSz2YK9aWZkF7uwhW1xO/WTdJcDH2i0VV1+E62s
bZYVxe6z5Ry2ga618jPz7LDGxJrne06p7uXNOil1P39RImUGzI5hddDja29I3SeWRwECDJVSOZRh
BO+Yk5BdHmuSwq+R7kXL2iijAbsrbzhdoKKQVBxraUywB7R6zJts0jFp9xRJJoIQMzISJvJsq5BU
p7orZP3kd0Zmub8AmRQ8bu/shf5znITj/6xTRq6H36BPG/kt3rHBW26JEM5P2kicynGM2g0iIt68
rMt2AqUPzs+h7hZDCWDLIe2hcvMQ13AxZItd4dIgU+QjLUtOxWDRqoub8ldpWU0tiwVIbQiFHHqZ
L2fFBYETmicITAFTjo5vq+iGDEzlKMp8JLzt0fkuheP7SgfZ/AEm1z9xOJAJzUd2fZe9Jss5RCRs
T+A8vaqWuqs0TnYER//03kJ45xnEK1GF8QB237SXhxLHMh9ZnuIscEELpJvo51xqvNwWhZw6i4/1
hXBdMGxTXjCOg2+t/hMy4Cum2iT1dAU1s5Z4ESB8/azifWUXvAkswWZtO7zpZuUeAEbxiE1NJyfs
HNAOxqAdk9rvED45bQ+VhcrzPtiC6Qopy+iDX/oIwGnGsWDQYYzNDphXKR914v63e9tbASqni/Jr
ppEB/W3LFfTXlAaQfQlBSU8n5oP5llJQ0BLnweXFbFrS7xjH4ipmKkp5y8LKJCYAhQBSwsmRpnbe
wEukru2ur87rDlq/3jdj8wj14ibbefAaq2pY+pfDBnYo9oElyHjLynE5GG8fnDrcdDLWpy17rA2y
JxXf7zwmZ1ki/NfBNETh12YunVR1pKK9aTxMNvIfxYeATPZ0JueXz0YdUfUjtKdyZk19ptTFi5RK
qqxMaTSvCvSL9F9NNeSz9c+9rGsr3xd4qI/p2YlcICgdoY+QtzARJ0EagFeBby9VtNYpxHqcT2Ib
DHzk2A2d1mEbvqNCkcSl2DRI83SRCQnNwSPqSdYWORTY329+UUA8MIErRmtwWy90gz99mgrZKBam
e5henlsYu84s01QusZWTe3mRRXTUTYQD9HrQNjn5ERUVBrsz1KJFZ6Pj/kRUWqJ1sERaOzd7GGhq
ijXAsZpKjBTRRiL0MwwE9Tz6DYYEibNjdgHCABQoe2PhV0qSFLfKLIc+KZrF9J6IYZjxehqQdllJ
0eIiMmzwaIeSdlGOHL/NCnbu4K1kDOqH0FHM8FU7GhNWInk5H15f6EZ5YpXWWBs8mHcxy4NXwacr
88Iq9oUzk4Vc7yVX4fYANP6HYfORY0GjI4j7cE3RPB69exz2+mxDpSCJu2iZyoC3q2mUYd/tIazx
GsmyuHE/81Xr4BE1tmDsCYkzTtT6bcwdBjULo2ExBegDrntvA8doqa+EGbt4ZeeT1fa4b8wU9v8u
O8sg6uovprJH4JEtITEoB7qpAuMtRh71pLDQFAOO6HKbHbdL8WNeFC4V4M23MW55cm87vqfE97xL
cZju6JnjTgs+evTJmDy6HXGfj3/lQCg8Hnov5PjPvJ5Y1LNqrE1Y7UeuC/pUWrzsUmvM22yk83i7
6cp74rxj4dn5sT27fZLEfUvARz+ur2faZ1WHW01VkyOahKGxpcTwZCTa4C0n3ifL+BrYUNar3dn5
aK7Fw7Z8vQA8dVoOCdFI4cpD/nl0D8Lc7XZ4T/nNDiNSy1Z4Z7ipZGv+w1hf9E6tFpiNSvNIVlwC
uZ1bz4w1+hMz0n/qVvBiA8V9K66+rPDqF/K9Djki6DQDgMuS3ppzBZLvHZXuTBiZ99X8vmD3ahNV
aDzMEXCCsiMiHMBnoJiNcYyqqrVI9KYIKaFUXCLsTgh9r7v7jwS0qYT+GgfaNi92ocCCILz3j6fN
Xe75V0ayMYKkUW16gxfRYVZuXJFxzbdPJX9TiM1CodIvhKNbkEe3lTFsuQ9f2KAfErbKvF6IrPuK
bLcYbv1Z7ZEQeWQt/poLWPVtnnJrI9wGaNLYX7/aVMSkQjW+HgyoUL/UYOdFU+Hsj3t6HzwXsjBf
8eH4ToVyoXkGDX4hELBSYCsOBmWNKMAuxJaZIotIX6jbESe+WgMrDCGP33COkEfj62HiTiQSol7f
WrNmo6X1OB5fCy0PDqgiNEKNuL0qXGZg3OiQaD/jliGGDhLVMampZp2HX+AiMG1vmuKVdBTohGcy
MlPMQJQRP/o+cVOzN+AJxN8JsRfbcftqFNl9xFhNSGl28TEM7QV3KXrsLg/Lm7AlMjCptOXqpgd2
KMDOyVUQ2ZBukJvj8VI9MSGVtSaRBVnFYAGHSBY0OM/AB+zZA4v6bE+EsPRoDOHxSxAtU+BV+GFC
JkMbjrk+ag1VXsmcYiw2L+F5TgYT7+RIeUZhNNfJhns0MWYUMRcqlRFt3Jl0QlCSlPWTcZhLLMDI
4ZLVoMAZBGFBxu/ILtN1jTzTO2jlOZQMlLAC4DGHSUaC14LGCberRvB7gRn7H4BXNwpcphG9hpYh
i0hNrxj5dShVERwep+8FebAKQRYrns17H1MsLMASXkQVqC6Rrl228l53pgokz8WTSLdta8dN0hSG
dCIOixsF/lyIqeKSy6BxJ2XspEzRSmy9pq/BBRWsRX62ul7TMMq3ITlICruqJihhpAnKV7FMKPjs
HJ1eaKrLmtdqqCqdz/qCEDB/1o5tzgxYiV7eM+GAaWdPUO7Du9ecg6n7nu4sn0eOR2lPB+I3Cd+v
fTiiPhM/2EgX8Lsdzw1DdhclD7Nqa3xYqpHm4Xgi1VbQwBc9dF/Uo0rawaZzxL0gOMSCYp8APTMs
uXEu63Ym89TZKNFG1hj+/IqfW48m/hE7Z+dQNWaqm4Ab9rNjuhjqFuDYJ7YVE/J2vr8rxIe+r7Cp
TcOjc40dFHY9zGglByBLyRAQ7hNDHM1xh9tEqLnRqXowO0CrUEMr6lqTPhFU60Lc+E6AN60vrAWF
Ld0w9uGq/7tYGrwA6SOg2wmJGXlvZgntIBKZtGsSe9yUBWa4V78Q7Oa6ReJBEnbvh8NDkMPRgRyN
hyFHAxS84/hCiBQ/Kzh2I5/9KkOG9HozW5ihgqBNH0sdS5Yw8zbAphHcP57NRr3N1BVL61NyfZM/
/25YLzJrzmixiGir5/OgRDfWqG7pwbrsoPMPlwWbAqc1zXIoARk3L0+4kmQ3T0WLYxu2uYzHDn0/
U0o9LAZl6wAxY4WVeaGh+WbDqNJ0zTpJoqaieVYhGe+PQbWwq6r2eSgZChcIh0dnPh5+HGmH0UdC
bUTWegRtAiOMtfsszuOYfX8EioxJkZxUh5OZuxP4h7VQ2x1brAClyRiqcMJJWF+epSYnX3sCKC/y
3GfP+PbzigNjsLSNS9vEGs9lgNVtam4+DZsOWY1zT7XMYTgAZnp9PYvuFhpSfE0+O58WKfuNMV0Y
wl/do+H0qdBEqIPbzTMpMcRAxG92e3XZlPVf/PC80aC0uh+arxufR3xdoyDU5vDi8e2FjPjgd9mc
8IyJMkIe1EATedxE1/piAWvEAo+FjxZuIO7B849iju32DlTgXgoPcc5n9yAGgZ0p17PK0FVt5m+N
ApFR5tnPwL/wptahU0qAIT6XPvdyy2hl00JpF+59MY1rRSUtk0AbWVyN3+P6zj/lLnENI1mnPWoE
nXaoHsTQdL9ejp1ckw8R8YUBAh1SEJOQ49+E9d/5gZaWt+7q3pwQ8rF/OI23zWQ4LH1GvewlQr63
E3Ab+70x/8pV/B3KVeaJcJDQ5HfMaFDQWvK+rPnejmRnQGw9KkwodBtbwfpTOZ8NyvbYSlWycWYX
yWKzZC/+gQgvsh4K+Xw0e/bRrpJvDVYvHahKDbf1U687NNAX+6YrdyYsEHia9pWAH9aHdU74JYV1
yTFEkl+J0pH8mWXrRY3ShfjX5+P/zsZRhR4RAWnRZ0IyupzVp8L8HcDILL/Phb4T+F8+J6P/JLEX
MW5EJSZsdI5dl8fospXC2YY6lOE8nrU/QFSkXHQOkuBu/N1GegPvhaue76amQBu65jbhWnRZF3Vw
TGqr4Nmoc/Vml9zb/IWQn41LIvni+92M1R81nf3O/Vp28iOVgLfOTkEHJduNnByDdbE7IR0K9iMX
9Nk93zebkpYPoTa+iFRw5rIu7VWllI0FBa07tY0DV1R29cb3/WRYA3+oooghnjGyJzlkB1QeZXfX
OF8/QmJYNG1VskMTXPEWZdfgm+wgfTJS1pkaT6vG9YYaJJ6mWZHjkiY6qyWt2ekv+VxlbjoI37VL
kj/wIF+1ind3Pgg3zCBaHyYg2p39AT5dvUIa6uqBBL5VqKw17u3xJt+P/phlCcKtxc4TW09RHFJe
NohJnL/dApxzxQmZJrTXP9iS5I0Z4NRGDVcD8hBBCU5Tx8e/tzC4iLA8EyaSwFJTzMaLSFexHQ1r
RdHcNUHCVGE3pg1DSvLBqkZnVCQb/Pn08T6UQhx/1rZTLMoVU1+atdqFgKoevhf/6xL/mEkJwzmi
OyvIs5jPzdGQwbzS2ZJJuyQx6wNZvuWKnRI19IjcOqdeEma6W4ZV09NRHOd11E83C3pJYVYWevvn
fx8igsVicFWtcS/yNkHptYEeAD3qTzmrG1CNmpnTKJ5KfE4WyopVv4qPEBVyDeZsOUT3imocHyrK
jDUMCkY6r3OF13XrJZCEXZ0/K6Hh8yTnnDkbkqlDCVRwvzaAw+JuKO0AB6A4JoFVKCP4jgbgcP+t
3u6tO+xVhkY65JEbRq8vZ6DjCH58T7GsYV3goK+VWAlv6KEToSjugLEi/7T2jPlLxdbpZjalV4qg
tI1oF3GJPmT2bgS+hoKcj9qeRD3gEEY+dSddS2kSnPAyRj/bLazdiU4yFB3lDQsSx975nvRa7olE
ZLkm2qUqfHz+teAeVOQCdSlu1ISPKaCb6YwTU0CFstiQSs4ad4Or4P95M4wK+vlPEafkCOSgnJW9
S8NY54snxEpS2FA/bR3zMRRlrJ3OUz+6NrQ3iXXqY4nPqZSMeDLw/jHR+78EMrZ/JT4TWnskGHJ3
UG+Nyb+huAl4I2oKp9LqOwBU7xGLk1rjzklsKZktahUoVreKlbunUevvoZzQbZpe1zd+blePqeiE
+u12Q+JhD0ju2+uihgy+Zy7ck5RYqV9Ej0JSehSQDcEnAqk10+JQ0TZQnJ2j89VUrPi7Q1Co6FMW
aoKLhOQ6rmuhWmAtgQtC+JhgbFAqRkyezLoE2gxOLDNDzxClxy/ZC8AZVyM19Uo2AsAYneAmcbfS
5Vs3Ytq4wR2nmS5BJ9ESkAoWCGl0vAOdCXquQNg8rGhThA6OelE4zqeJlGgzAQasl8nIh/GiHB9i
dHkCq4e8FQiXrnYn2ac0NHysuoMYOmEH8XBfMB8iD4fLTo2xmGtqvSdMolWtA79PXD27wKnvaPvt
Zq3KkZZFnqZ2uPaib9PhLgw6P25Wtzp2g2leDZHyX9U4DgwpxggRvXZFPFbMkQuU5b69s/Yqbr+m
W0adaSDnIqw+w0AQ8MhEoRp/jjE/q8hikZF+apswSIc1FzW72b4HzQIoc/D5YkrcNhAXL6XUlJps
VCUEFbon+MPX41ExyMJ/v9894nvrqGchkccBslu36PSru1k0qFyq58CGjeIYfzkmJf8J4PKkaK8D
iEte9AEHOCLBq5wA49B/EiaAICazAUtzZNY/MCZhHI/+XOZk1HIXs4RQ/qDAPJBHLVcqInMeovJr
hNpUoGkt42F2hfhfPXlP0LQNea1XlMakyXoRHuTca1R727pfpBgriNbFYWZofIFoZznId9fnLlxO
N1E4iT79/pJUAT5d41u/HrbmTY66MRKMgG2C8fsZo8jQzwdd7nmdBTpVoT8Tmbq4D1aDmCkjhzfF
wY3SvZVWWm1rx/GkZBG3jRCrwQIs8vPyssPaZvPZqA4C12GMy54eH4MOKo5Rmf5Nu9XPAFg593J8
PCLcVbEVMbus2jAsSfEmKjUQvi8kI5AP7nhjBlJ2srhryUNW73C1hWF6SrTdZlKjc4S9CGCZSGmn
/DCKqHVWYcFwAgr/Uum4Z1J9HYO0cu4PzILkpHoRYq2KUvNJmjH6BKCwBfvUJBTxDKhB/cqSRmUz
sAacMJ3fT3KJzDyg6ZZrGybAq5GhxXb0iYqkd4yZp4zwfzin3p8B12j1KzoLqSj+3wq9HTfoqtUf
LUHEAFVswja8x3FgL9s9KX8loCLvHSZdlh5MzUJZDKuDa8XABHLL3tKQWztK73LnZYWtK3/U5wjp
MTtGLq+KcnrHuYCR+Jsr2HphkbRnRn7GdBS4j+tA8bxNKYvdGrwRS//smc3AM3+zEzZPyVvUUlXV
pFKfgw4Cm919+WO8PlG3DctjAfG3YCee6/cm4aN2DkEKFR+89/BpBN6heVktWVKW8JSd/YRAELW9
m18pGMVoWD36XBffsMAFAvQ0FJesrXAGJCP4JnxPT57YM5LVTokOsnMgjE2ev2NDr2u3BY0y/hAv
zyOqGdGE0EBJ3pzHDuujk6QidTO6pwvRAQtYnwnMikBel3vf5oAE5FeEVOH5uJ5UtTyvon1jqxQ9
jiB+m0pf93yCpM1Y+SXaqsQPzcPXCCJvIwblpAcIk+AEMX4W9YbrpENBQjcGfxmYLgj7USHBbsnx
/VxQeZAAoB5tn6/h9N14Q7a5a/DtY3CafAP01nU+FV+yeO1GpIPfV3tRSO1r9IJ6aP/owBOoAcH0
Tlksu7scX1At5yXzwggQL/X5lAfgEN3W7gJUvmBIKcacLjZuWX6qrJFgguWLUkp4nGbJMWOILByQ
NcnCklGTjstv9c6ez+UEzya7fAYLGrSBV1Jcij0oAJE3Y27Yv5VM5NahQnK4nRO5XUL4Shgpy3KY
Es/HRyvqjVIZSkObp/jGmDOjeIvj+8eD0N3ie5RUP2agdo97KM1++2mmKsoK9CzufQdYX0tSP2WP
jpY1aI/qJOs92u/YN6X3CRbKMW0m9+COSkQ0v4zW7QroKOeCsIr46jk8iycW0GK1tdqXXzV4/ohZ
Lh3793WbMwp80M1s1RTspjZSjwvV4aL2RcX8iA7s7ai5s6dq9PCIxdWLyAD8eABk/Uyqrwg0NJUv
ja4iPLqceliWSZMDWNMa+tAFDt1UM9smbD9VM7nh6UOCVD8VUwkP+GbVBaCyF+9FKwpCKXqqqpBu
mV/5XLe2r0rei9XM6zBZtKS+R87Ro2kbwGIJ5xyUZ65X+Bko6qSyvBaL9cK4plvJ6GyysIvCi8u8
Zcq1hHu+LYqbqn8B0Y5wkDMRseIrIl9VlB1cjOiKh1Pfl7s5OjnRCgve4QEBF9frdXSKEpcFvwzd
gzhBdcu6z+f4zKqxtWFzhqXqc0yYFTMlz4Jvg6nIKJdTT9jafvj8Na77RzjRDzR9gAW2N5JDX0E2
D9cuuR8sODTTvQDBFCmvPd9VQJOvXW+7lOeRaG/kCvfY1ISt0Js3uxTDHbxR31LnBlGofHnExXNL
zXlkDilhpLQYYTdTJZIfCn9hFXf7a9lctVEG5SmudxRrVoR4Ibu41LOMMtc7m32l8JkS8NFuewnZ
EDXZYf/4qsTyncRUETS/AbmtySD/NbL17vSsesETsHlK/iDn1JZgyyXKkyM4jkPhHAm4Gz89vmUR
eRAwbOIH03X5eJUfq0HPhsrEqQ9eA+Ou1MGre8gVStByWadEffcl5g30Iw6h4wqJvsCoZAf+bPri
MqQ5pdYwMh1wWL9O7TtcGzkHShK8g6No8AFc4VbMmHL/Pmqy1Y/eWCiSd0WHYcpa1ltRi+lItj/6
HiHww7f4cQh0syawWCrDf24dtjBIkAZWXDGH5P5WcHigUeZTsaeo35Hhl2IAL4RN60PpbIIqEGE6
EK1J1ua6dnW//pBA7TYsSQDP3Us2yYJRk5KMuvAZnGKurMk9q+bQJsHViHBG+VtdEXGvrACjLNW2
SaJGh5ozopbM8SfReP+0VHl/8hv9b6DWO7YLMTBYvfpxLUUievfIOQkIGmXBLOrYGlkfh8FpAjLO
pb3q0UMv/sH+oMz/hWo1PWQ7qvCjEZF42rw6yZjaK4H8RexLfEiD90BhMC9pINgzgTmMTbGLaDBt
gx/JJ1+2Reg0Fz6N9DIe8RizJSSn+ro6oOGFpT+A0G2cCghhQNokOtWFyUP0A07LWR4jX6Zoqn1v
XHiBSgmA4hcRUEIYwpnNI1ZNqCF/hvzvIvQsHmsqPXwCmZmxCD2jD5csM9CsYmLYIzYl+fsQFKmZ
ebK3DkJWJLnQsifszpzdSX/NQuhd/sJpMegG7FY79cGT+ng16qD/2G6v1pGkOWy9qhvf9ozz41Ky
4NkeKd3Jga+gZDl5TDCA2gpxznVz+UVaYj7R7ZH6Z68H+1QkWjdR7Uof0g3DjAFan8o8iisaVdXF
hzYYlvOrmmLeYTKkxZ6FEsvTT32ZzwNqVBW9+cwkPR7MYX/k2dIaNl2hAd9pbXuCdApiH000Obn2
/0IPaZZ++dM+XbYJ9oqhRmeu2IZe9//ZaFGQaVaX1hV2ctptHvlSCNFZaZpKDFO6bNR2dHdocPvQ
vyFsXD6rqx5IplDDgBQo9lcPhqPq+ef45kXIDYUdLhXrTF/B/MZGxbwNRplmpscP2jPezcwaV0NR
deHJU5vGCsauSxcpS4NkmI7xbdsPL6pMHW2sxMCb253VggnM69jq6Q4xAB1a6HLnqZAf1RPkOB4C
vSRQ+UlC9E/KuHRtH9f92W7lUr0koFfWCpM9gfbTbJbMjegmTSHEl021zUMbeucLzIeu3x7NhonQ
49YaaFoBZK1MEmSldv079SBoHbHR9xX8+4xRAlNA4vVputG2pys5S5bbJlYJjfyseJkYjvnyaeSn
j6PD41MAs8MABr02BylaXIudHEvYNTnGspYk8DGan0EERRCgYD3oVzSgLJxXxLSnUf8MHmb42OhC
G3su9OdYcAnCCi5zqLjFSnv01bQgwlOqOAuUlNXcuRMN0kp87j1mPGDAeTSPci9ktUioXOQdDbGq
kPTKjQCqY+xtp+DSXe8XOywM6pbkbIMcBqKiM4ALHSPEjeM6PhMOPUgMvbsO+ddJF0A6078DhJxv
yZ7U2Kc0ykz5ihbbsoVZTnLNgG5eLrM7d3dhVL+mu0DGsKdXElwMurmDI+KGPwuuhoLjpCFKTmv4
+bpRFabaTKRysrESMIqbaQtha9y8QIKS1GHQTDnb/HmdOxtKon/DnEfaPPAM+8yb/FRZ8Z/KOLsk
ijJQuF9bXhqoSWJLHMeeqQvqr5uegyP/Muj3lsFPI2umL7Sqps1/W+4DcHagFJvwLsFqq2xcbSdg
VTuSlT5oaG8s30ljz2Bxy/jBsDtXdAaR0+kAxNe0zL3drL62Np8gn0fpfs1rjx8sVFKqSYcznlXk
aJqLCkTBA6Edt0e/4tNDryGbPlu82lg68TLHzzP4vX+Ki6/T3bCPj9POt8nqs3qu0wO5/so7nVhS
EjAPx5iqgxlQGOSchPBDkjqoYN3TwMdu6Scun8HxtDEhoeZIiW5MfwcfbcuiNUAbvOlZzQNGT5Vw
XAfOYuEp1QcFCNPcnD6jjuq+DXfctvp+KxRfZgk2kZaUcSFey6anhS/YwmPrGY8E0GaLlTdfwI8A
6YJc3ToCgrgO7yY/H4dECZ9bBOoTLP/LooS4A7WJNj17vn92gFEJBMZDCPNoJqZcofutCZuZ4Omf
/88lXztx9lQS2xSx4IRMFqAP0bYiStdnMzk2Fxm6qzK+dos9CU+HHd4vv9V6zZhikffzxpsix6y3
oM5fGHL6bZ73LJGoPwLcc+JWM30m2Z/Dw+AG8LV5aHuId40ktQkAMHFN5buvzBkCC4JiG8h7udfl
WWgjwvGcGUYdSbvtRt1NDi6rTzWKRX6WOnzKVp+/8+YlLb9A5jBXT5Yz8pONPoCDXPm+KPTEUzcY
NX/SQO/ACYPCkrXiaIh5bUQa/9OWpNGeN/9j8KBOCQ7fSPpztb7nNBcsq6aS0diaaGFW+AuH72XJ
xKYPX3YjtY3kGqEmB+HDEZgRJUeWhV67DisiET9ADC1Neeuj7l9cYLIG8v28AkuHl7DTmPsQjPC4
3bexJtq4ODidB03PJOtjOSqpxGcNI4xh4+h6CA3SPEOI43VIH7p8LFUc6ZZ+T5zCCXND2bLmpEpi
ksaozRq+Md05dS2RATWULYMRRYIJuBE+tukYI0XE9H5xdXs3A4592lluZ2f0kodR2LiZgTXaNzNe
YrgkG5nlv7NRdXstgRiylQgikdBu1xDXCPhtV7gNDl0WJ0kdQfqFHinCrS80bESxjuTWTF8V7er6
YZmXmSMsjiKt7Dzn1HQ+yvhyotJ+FUzGdPapDo/rLJ+DLoz19b2J2J6zNOE/cwnOsB1Y9+zHZvsb
qIeb6t7bxZ4vzTO9vkyXlGrXy9J8ZqmSs+uPdmKBNTJHeB+bHwx2QjMF+UXbHwaRww62ReQi/Q8M
2nlceW5GoHA2SJdww3bgfdEIDyT9j1b4lY5X5juO0uOWDBfHQ0YXMyl3+LOh82oEteSHrVXruaeT
JBCaI6KBU5o3+vwoCwMCJl4rnlRJ4PRRUqozbq4ScTeuwnPeC3R06xee4WgSStrL5fPQjpaknidO
VMfa9l50BZ3/ImBsCzKDfn82WHOkwRW5tLrDBd2r3EvDyVdznndEAq1l8Olkvl84OVwiZDeBkECX
ELH6tigoiQ+busMIEcFOLM77BZWi9BFJ5beLKUjv151inL2rJHvyOIzR5KiqShkxJ10ojoGSUyM9
QZWDkpv9FrUJeL0PeKQHOaIaJxH2PjO/6k55It6nAM65XjzKWCiRVXBlszvPAgwtMQyGLhMC3BCi
zfKzyVSxQ5W4L23ZJ64iC5wVw4lSdjJvpxsBJM8dmUDNs+0RI5tCHJ+AsNknIhBcWBUETKNCLK59
bestAvOHNYjNQASZiYXdrA1L2+/juEz1gxXCtxqZU9xYYzSKq04HjKX4eEvGboEGxGYEW9vuXLxU
aChwy9BxDWxSSETiNZPSooDK7Y4xTXHBZehrsi5gpQ+K+zRS8e6wd4iABMlYQ/ysNoYq/yzMi/wN
u2SPFYudN6ms8Ccd95tVsA0b3UZUdWAjGiHfN2vkCTMWzYa9h3w+qs6BlBFNEyxWsJoREJ5sdSUN
AaCKcN6cccYzOlLA7c7xzlcNwQt2Xv96ive4bWssWemvqwRdLpvJCpf+0GCe0aqxf437k28PWWFF
rI9cSOEYcZgSQ+bR7CrjM22qE6k6mtobV3Wiaovh/wqd31KxIo49DDb/nkuXlmYqBQmcNFDXNp00
BJfgUpjp4MT4aPZ/CcoYM/h8stDqh5nMOQ2wbNr9UEG/mfhHPtPbFH/8dXdMceU3wOr/qNIH+84+
AZ8i3uhpm22TIQp/JbCMKkslFjoIhC/EOj/6qkvLDLBZG7cyJEWSIz3Uhlfdgv9stERT28X79Za8
fPgQPEmH+/r3aQiPKWH/pT+IM6qpCQJ3iFZxCSRj3qooWf/OKosiJcZsxp3TB6FeKWLM4yooTw3H
9oNiviBGQA9jDUJMVZ2BD0Htub051Iizlfhwj6wGu/4oOobjDJFOy5kmjgUnhwi+i+KLhpuaEE02
Y4cXHehpcGUSs2PbQoNK+WoUYXkvKL1V+VcKfRM7wu0YXb72PZwauaJgxxX9uBqzaRv2Pr8kvxtm
zLVUhJ/vFt0xAS3talrH0+1QQafg3aXl+gMNPr0cIUgeOh2dxjTtTcKt9y/SYFPKrIeRYAf/WhuO
1z5rd3A1ZNZXrc7Tfi3cMrFx4YR61AKO0z0WZuV9jmD2DLK1zmHD1PYncj1oJQijQxd7eMjR1nIu
Au9GbbMCTZ9L4aTmbMgy9k3kwJpgh4PkYWVvkfXGA08jQwTVfEh+xLAVRtjysYyHM4dh8cUMF2Pn
jD0xptB8ODeO5wGHMeu0jEf8fNJHqWsZH2toOZ2ioPjEpaNCf0+h7b7jSQkx281T8agCuZ3puwEw
y5TNQdj3ynvsuXpJXWQ3sAQ3dZxPhA3vGkn8+Xm84POWG79YW4VNU9QAz2lVM22mZ2dnYdOM1aBF
eMkjieOYqoVbchFiVZgucoKFI7vjwD9ZWIGRof9r+WMwlrUbyGn6W1isFc+eVSTbRyePeUBlYdR/
pxtRdvnUxUpHuPaDq7mdujdmRfnVMElMP+g9jOaTHjukKmRHd8VLkwfpvSDENFiiNykv5oMCMC/D
GCQMpDZf9YjVFKaZxxvNeGPU5i8qIFAoybGKK4/Q1Y/UF+BdWKH9ISGKoUVhYRSTHJloNLeMbSl0
0C6M1jFC3zCOtUvFyaap5vGBR+iIQ5Y7PGv5hJ02NVJ05pKvLMBzdYAzzJP4EiGZ9B9g9voiR902
6me60iF7ct5AuMT0/wX6RXTsMbasToteL/7NA+XiHEHBnv4OBQEsX5r5IEvNFo1fM+EhcVwR7EsI
lHshantUZG6CbWTZ9gvWDGNX33J1i7iN1b0cQGCcy5mOqK3kKY0kotIHOX1LtixvBcRa8GWwpekW
9L1k9NGRWPpr7cGEi7syOPleZXEZlvOxE+nkr4+mt1JgdAfrIKCq/eA3Hj7NwzJJ3pWhvdlCN6YK
08AyQCp9vrkzxQFrhxvnALUzUYSDivUfdXFLSIwXtQm0pgLRBmUmVFm+LTd/IQxo2VljXeLCBJYJ
XRquKvbT8shNJNRrB36YRD9MARcMhD63JUmoWqFgL6GQIkCRtqRcZKKsXTX2HcgjvTBZ0m5X4dWQ
SUZ47+oL9wkwUH63H0/1GMhRvJu9fqgzLJTKVxOQ+WTNT1mgAinhiC0PlyO+01HFHuAohYz3SzPP
IC3rCFGX/BAWuGfoJmGh9CX2z0bPTTP3j/wRBjgTC8t35XXJ05RllxpyRzqjqLhlf6Rgan6F79xj
KQqrT2JFyJ2ycI6ayLwgEZcBFGacuRGVOb7EO/mOKi0bWJJotUg84r6TbEmkpeWk88VKj5Fp8Yn2
Jl6JfsN04vzygadLyzyV3UNxplLpnDulpUD6tKQ1S7juuQIIznkScFhcd8K5CsxWnhDPi3jiOQF8
7FbWX3MTKSu+erhl8L9gi1Fe6cGRwbKdfEYgEVF2atAvc90amn/Dz70pryNuPFuZfxmxekJcfpWQ
LjOraqyriUqY1NeTsIF2IrH3Q1IBGLfF8+dbnRu1mCli4qZ3YXd2cob2zQQTCFNg20xSGpWucF7Y
r91B3W0E5Ez19zkE4zZrKHOSZQ48c4QNFV+CMwQWxqJlusDZWuAaDBbbbwBTSYmUhe3zCUfw1Kqu
ewCaWXLwYpT/3eRW4WoXi/csG7k5NwHxuEBIMNH+EskGD2OY1pL0adDuLZBUaDIKtyqnEy89ncd7
8dOY9o7OB9MexVCCencp4yVF0NWgZbFkMYQhpFB6yFVW0cEur8ShowN5nUWeXzYK5YTe9MJuNhqZ
9hrFrldy8AWaLDQUH1H6ZftcIIENijbuB1LTGiXbBfcDyumTL5EWZB4/DPmhaYfCJQTtuBy2fsIx
ohXXYZZ7l+0NAuduI+ggq7dd9XRsNULb7Lf+i3JyY1dsz9z9YQBWobZP/FRHUtXKYgsIbgoRSElB
WPCi2r0O7wCt7ZA3G5DN/EM+4EjdY9FIjNyCMswa5FfAphxTQEP/tc7moj6tU+ete5mn+Z9CRggc
wKOp+FUH+YzBMdlvD36TLa3js/8qfreah8lHNZQKTastfjj6SgOIfSHCYEKx8HnsDVx+scFSYWml
lvWH7PO/rDWfHLUat1lfS1U44xJ2Fog0dAYaJoBPuGGhYTZq+E9rQ/2IgcGh1Wu5GhKdHBUyqnBI
+3p2JR2qePr7m0rV4UZIPgNV5j5BezQdkULUIhtY5LUOTIlG6V9PmR5WIw+qdCegM8sfQHXi2UpH
BDVU8vs5MwDs3MeD8Zjt3mV0qQkufJ/r5bGoorv/q5Heget2a/gyUqVFZsbZEu85/xVzw1/t5QlM
mzeVxPu/BRUQDQ7lnNAFoVlp2iAYWziqh0EeyqucQnzY0Mm8s56DE1pimcFzLFT5UDhPOJahpBJH
DxL4l15DgYwS1k3vNbMJ8Pjcihm3Msn7ECnt/o8lL7QywP28qRG9UV2FrP4stwyiR+IlEepmhiXM
h7A5//0E5Dhg0yb4cCp5lKZ17t/BuPi2F1/vAfmUrE2rTfgIl75VcMK2t3MKfq3HZqWzZpMW3dou
+dR33TqMoRbQf5wBAFsmPfHAAno3PlzvSA0rPvy+spshGXjH2QQVgPyZ4xGSEqM1edQIi5GXkyLM
Kvu84YZeCjAiYmBsgikm2KIazQjqkKZcgex57adebOGauAZ7JRnJELi3DpXOqJWxI/TYMu3ZJQeI
hnh1XYY4Tc1efT/0WYdUhAv8OslTQ8BJ8XeyvgFBamEeTRP5SdRfykSH48O43cXYMPPk3pwvXrX8
4EJnCnmfSFz2P2/Qc15s4B7gJKJDFnT0ApHiy/16bV9tkYPOTzhuuMlOOGP+CG3TOG1kgnKYx7Qu
MKpKG05BJ5T0NQIH/eIzBxxTCAfqoinj7sVnd02+V5x70jTrJGKEyKneDmbSj7M1xoDU8REH6yML
WPEAkg3ssFPt8be8TYopZFbNVpiuLWbsS4PPUU7T5rrkvG3uo9yn92YbmPfsTavicfO5C3TMBnyA
RXuQ2IxlUXVw993Vvr7l6P8zzNUA69QQm2hAmc8181fPXDNYTGBkMa6kSJdR3c/vDMl2C0NKAjQX
e7lDEFyXdeAmCpgLW0iaugfl4t3SFEXKssi8F0EeJJGTpGufEa0g754Lj/dUnId7H8etsHkiLWcY
3x8H3hUJHsYf96h0W9BbihjY0qmahITTKqvUGmC5rcuAJMwID7a7BaS0LbKjlH64VtrtVyu+Ol0s
hNRek2TuVlzsoTgouecpYpQY42MjYZ73XUHmw8gr5yVjXLq+uX/I5eygoeu5i7tLa461+4sqAMCc
TKEgLOr1Nxr1GqlwHGhZnIIZIQ8cGJ2X0Q2tQBQ/c/C1jsCwAyDsnys+hrJuiOLz7AWxfyB4/nOj
Q2mzAVln0LJ5fvmP2kNjIrMMj1tZqtrvQcULDn5VZSjNYvpCqxy93I8ia6Biuhz1gXQJnpRgE/4y
d1YhHzTmSPXbqJpqGYhXyR5v5m3Q7fiVYikTyWlGx1uHsu9XfU1kx3lI8de73C7wuecX2a8+sKG0
hqQPxsahf3annnfT0AkfZPlJCeEeO2JMPjXTdkuKn33h6uk5jiIbnc8N9nFrQxGzeo0OlJldjPc0
qZxzxHn8xte+fJHn22fPHZV50g70aPJp0ueVcQLzFEPbHDqBsuliOh2BEJwf2pHOrW1fKZhdnV2J
3JJ93NuRcH7KDkIXKXBjNK7oKov6JPDPp8hm8b0QRoFhltG6YT39D16tfd3efZHmx8gV9LekghUa
33Ov1LAXqfGhxDjd+u9sLck+flzd3lE991kgPzduxEVRImEVxnWP3aTM/3cKJMAuxqxChqe8VI7c
zjHrAUSCOtRf0P73l4ACtU3YqClDlRiH0cgSr3dxkJpCojGohsaHC/kRMu6Kp5gjrvd8RFiXP+nC
2hmE2S7oQwgy7p/wdPxDpNz3o3c/0Nm7g5XNAG9Ho3jnbdm/khLpb9ZfQwxcZ/FXdZ96RO9gibyz
3I8Bjf8bw3iuMLcTJl+NLAPpezsFNDgkxrxhfFHohh9yecfop7Vf2bnDb/WpdZmEWzMChEw2bLOc
R+VHprbxXCy8rxdfmLYvphFq9zZvdTzQXqeH7ETsTFbQ4odtiT8xmCDs0DMnimgCLjZK9WxxHSK0
TKIPa8mbAZ+2Ez5q5cYfC3YgjrXphdjBEHUp/ixR7+xcdUZu/b1MoW/8XVWjWLa4EX2cdvsVSCij
4CXRHj9rHe7Fq+X/c6S++ExDQ712be8fOfMewCmEv9gDyKcSRsbmU2ajTVymO+0QvAUnE1XWKkZO
O8//PRd93g9iIAmwi5WCphtKq0PejqVC8N2LsO920XmqldjFqkOJ3S0ddtKz5LKb64yoPU7HCP2u
PNiR1PNcRs5cYPoQ4If7QGpFzWppPJaZ6TAh2mgJ+DrmNbeGVGMSJYQod4f5/j9bQpBK95KjNjo/
Wdo3hY+ump7S2Xks1X9McJCYponrAQW2E22KpDvM+Gae213CkZgXWOsi0LewX17d4/o5P64k81t9
OGYMmMTAn+tudto5KV5n06tYDwIjkad+rw1UvCw4n7tDUaiACYtd961HWhdouiWCWbFuTluBbrmo
NRSGDmINeK9/9J4e1wBfI95RFreffoDXshtz8s3u3x5duZGJRDXDnV/lhrqEHllC3oMgmk0VPioN
OkvZo2A4EVE0sy/HBFM+HMGa6emji1A12kZeTy6jmXh547h0w3U65GjzlZQdWqvT3jBcmYp71ZeJ
Dl71Jih5QRdcROSKEUh+HTEgjla3NtZOQYY2Tn4z7M240HGxRNZg0BAbT2vDwHjaJ6p9FYhecwLG
YKAxElYd31g3wX5WU4xuC/wxwRAOkRr1nWqkMUPO2emTPIhW5AHySI8qBPsB3WZe839DtRByuO62
kE6f4YmMDZeJ39JSbCxTnhQxBoHoKU1mCYKg35cr2yjJxp6iBrov8mQIDavv5Kugk/wUGYQ9WB78
4aSlWFg17Y1IvRw9ZuEJVnl/ndYySVYvjl1iWUOzsfSG90jPP6Ox4y9f7R2JyIG1QxRO9MLrqt6E
wFZ24qBiMsCJDlL/kOAYkvp3NRoNq9LTtRmFsIjlu0xSsoalrjBbjXX5vAESmechFZdhQDYMI8Az
F89ge6XynnzbyOolNODne0ElXKcNm97pZqIPYcHB5tzVnYgGrYXNJ3E4GmI5PBbRLslwF1aQWKWK
YxKzNmQ710miClKLiOQhLTBDJuDacAULWiZMbP4kfE3ZP5O44b1bDwIh+JrtM813ItSaB3iCZbPP
T5AO4kATWjsauy/zUsMB908MBoloE1fLs9tTAybz0lJ6toD15QIKLUCHWF4Bs9riNg2/XAi5I6zT
6beNKwnQVDbvHTmEbvQjhVy2JEMJFf5466h+Czz44s5jFCbcjs7UCklvyjBwjuQ+eqy3yCyCrjCp
ibrD9GgVyyu7rVJKNYmzQV8/gsTjF3f1437brRPW/KXdcXqILmba9TBqmzJ7seNq5AnxO/tbiIEM
5XeBlh8K0duRHUF/ffAc144f96HZiw3kPhOvREP8HysO5l+1MYH9JSSnb1w19RxE6qZQo+g0bJVE
86DwiYuqid2t+tuY1OchQudIWUwTCA4Zs63GCTt0oWglrLoOIXMym3/6Nn3ln1M33gZmbx2ZpSMb
i7noc7YkXS8rUKTagnGFrseRWzvgVnsQzMl+UtUTohivlZjoMtjp0Z6wgxgoeOieFumDsLmTsGIt
DuuPYJ2kHo5v7/JFDpezF+NXZR9+GtYrln0x42YOhWfAey0dyHPHXmohqxY2HLE+lywd4HWDfetz
boK5MmN7lyD0ZhM/58yiyyzm0Sr168feq6QZzJbgDFZHqMxqFWJbqEP6UhWgiuvBA9sxbPsauIar
4jUYMidlMIvBdxTSfMou6/RYkwwgYcIc8s1++9qvDmrspEJYVOwA34iFxhaOYJ5uqS+rBOUVyJ4u
VXhR/XJmolVeh/LPCyDw9gT2oHAy6R8Y58zYSbGF0topgyBm9Dc3hWl8ofre0fX/agx5er3vEGo5
w57OODNv34W/x/ERvQchZE1MCOlT1oBvj/zC4W33HrczHmJORJRq6nj0Ng1Pe5WbFsnWZC6wf9eH
/tHTiBgcPgY0s9wMf7sfDwJHPobR4CLnh7qK/zih4ttF5BTZ5MNaghYH1t5KBanCu92ZQEAit1Bk
sLWGBAqIW+AtmodNkzm2PAcFYyxJp7oVxq1oyOf9pdRoUjVw68D32RT89UR3tz7/rmupB9gcwb/N
imwH9t5Q7GW0MuqhvK2G0m5vp+knSblmfguVC992D3GQSUt6PDdOoCdkfy5if0hHD2D2fRzCaCv/
IyiZVT0cYjJjUR1jpGcvlsQfmuvfCGDQL4enDlgnr19gZXg81ULq92GsCo5LIrtLtZUa5vykwVeS
P3w1gaQfntpF4f2NGHDxcArpzAM3I3optRLfGFdunNuLBF57uL7ihsb12WAj6AWP76KFbI3Pdwid
6P6Ivcvu1cQXPsfSZEkFJ1ZH3lod6hdqLYlE8ggSkI9WdEzbfQbo5Mu3rLEvErIvHrLFhaFU07Y+
F6kkjS3wQSt+M3CmRRz8+9Ryjm5jCXq+9p6u7jVqgeS7yqBICS56UVfDKbIphpOaIOY9LsKBgWq6
SzEx2aqp26a+fJRlAdodLGlh5Zmx+LkH8TCj6ZlZqxK0cXsenEVtx2Ao4GdmmOcZgTLHdp4Jdb7u
7b8QiHHrZkth2OoTzau+BlM7k4/MSmh3TNKqCkMpZLcNoQLUNZGjdtIplcS8cs4jxPf84/QN3uUE
qROgNCyYrX0loDaoafpAa2DKpqrBO2Oqn0G5bVGOthCT2efOjUuK9HAop3xgpcCYOB4/H4bOZBGR
vp1I7R30RuAT7jtb2RHg+IWdB1dlpfyfjPSig0bAP8aUbiQbY5vNN/lMDSkTK6dbZCb3Qwt7oFk4
KnXxSDfaBwwR2wJyTaVhiDCFVvSRtsQ+HcWU+e9Wahc47+zbgRvDKhFpxT8DqDYMZ0XfTF3dhzN2
tz0xzSKnZWeFW8iprwKWwSaIi9OszTf7bq59aO/LA0LOpn+F0Bmux4W3OXO0jtgQxsZxDLgLzThU
yyvuz1ToA9OE69gByij2n6PYlYf406aSFBA0CyCk/vmAQ9FENEugmn8PacnkOglzkDJ76E5QaL4x
bVVoAS4yThDvCjaPLjqbA+l7maAI5qu/uD1Ad2uO9JSsXRn+QIL9tdC23o0wQ/35qo2aEDnjLaOi
+WXKyCoGxEMUEMmGCcwSsiwVVK4Y+P5ozGMCTYc+7p2fVzk7IlH72v5zrPPDl0qrYy/Grs4+KiZU
xZcOvE9XgJade9t2b7BJXHdY0Ro+DD9feA2JRwWL+1sJrWV50oFB3nNnMgXLnkKtq7HyESatya3J
FuY1hy1oTgz/Fq0XuoERRruUU4QxAUCwfIlOrQANGblf6WVQ4SaqWCRvM+Y5F1OhYqHpQdpYTWG2
4Brb9TVB5FN8mEuqt6N7mLTNpS+8L+Z53s6u0RcS9+PkeuJ4hVEMM2SpjT/N3cuD5zbwx2v3HylY
1/PjbEz4ryw62tQzZOsconqqoOxZZc+k4+Vw0F78cxlXNTAzUcDRcKTTTGHKcQbFtpzyXVkT/XwR
wTRV3C0MJ7P72aIG46Yx9423MsnvUsYnthvJBTKDcfgJF4JwLVtdItV10LqgDD9O7YlCw8fnX3GD
UsJI4QNWhnn7n6YOUKfcG8Tsb72aKbMWR6Xan0OSYhIvEurjIwvciWf4rjxvW4xPbeXmVd8GkX4X
W9JTLycG9kS8kcE9ydZXKIT4d+Rdq8pnWHBWXMr/+gx9xKTHiuUJTXgz7BNKp5AHCEpLwsnVMWGb
NFfR9rXT1b2M+Q9E2/2R/17Z1MUTVUzCGFsFolBY6Q+18inmEVPxTivysw7RL2Xxaj/Yop9vYcrC
Bl03YazY04r+mJa4aK9h0ienBooEqKMHI2YNiBeaFj10Xc8P6gquyh18Uvus3QaRl0B6euliCjLz
MYywnOzAj2hEz1SkOhgcIdyiRBZodE/EvN91s6Q4R9ZsfTW+TEtm1tNSB1ql60u7cSo5xu/ukKei
2QCSqE2C7BQVm2K8nd4n+0Respmjzl+R+r6OJP2ALv9R0Nvt4JadTZwNTcwWttnxuODwIRsb9lw0
G33F+uG2eT18ZDCdLxpXv+DZRT+luLYQ5/BzWORFH8KSe2FJuOFm4ur3tvg5hiXdgDICON5qjVeU
0eBu6ZW2MToRBOL+rNkprgNiBlDImPk9Z9n0ybVnzhgbCvQd7xNfeEnvSYRKtd9/+ZdLgyYmbUx8
0d9Kbl3z/FFwE+3FBCgiKCYE5F++UjqxKjRmOsvRDJlGTYyH7+QOnCYDxe9WkAGTAUB9fLvlzqI2
7k5X/pO0szg+RREsDPr04FIVRdifQiAR2XVEBNe6S7c0KcdHpBtalkzpTVedmoKeBZhUCcNWaP1B
SoRxwuKEMRzfx5HDuZPvObRrfkbHeuxF01Tt79ILg4B1WjLifMsCW6oYKJiQSzQQ4AHPhYFgC6ix
ZYMM2jVJyjgjuCWel4TLMy0Qvd1z76iyE2FcblwEwp6wYhJE/OX0vJZRxYs2bU3asn7NFRbzUPRU
jPLFy9kwHx/xAyVJhhz1TWEtNmHmbGIX57QSMwVJRGu5u2Me2EW3hPkN+KsW0KzWTWf5ogwhvxf1
VMYioYHlHI1BvERSZO3Az8mjSAvUnDDGCMA18zKfg8Ismfoo5e2q+uNX8BNN9xd3+VXdeWFB0ibz
i12aTIj9O8Pm/sInHgirXLaKdF2wqEcQjKxeONfx5Gvt7QydnVnnZhwIFMtVEWw04L0DWfWGq+Iv
W6LDSclkXFdaYgv1OvoMajDiGHP/jNmcapYDFRTmYpL6h67M6VrnrVagtv5tYGmDhc/LFCoD+w5D
ftPPlM8ae6hz5u9joUS2dZiAhoyWhx6mzcEVbRExSwhTpXqzElb/rDz/FUpG2uW+W/7L1lHcMpIs
OKAiMlm4WkltT8qaRpkwdoQPX1x82Yy1Eu7vGNKawDrdbcBiuU+JCQEybN5p6RcDeKRqABBiSr2z
F4qP9Q+fmvGJQxbQHVP38LNbUfU3tgZlJWowtAITglwTAsbjprZRSL8EQ1CTcGW/RsWiMD1qNvMB
kSi/Qyzi7nTRZmJWLLh6cDc1FvdXFaAMMZGjVByKekydnVhrtFlQisB7awnv4aNqtJkP1wPTYU8F
82GqwF6pdNRp2e4ZnBhJ1q0YG5bbDhHBovNtt4RKv643yP/pMTzfX85EJ8rAj1PBWYDP4yFSrXsm
4sTs96xZThub0rHIbrpdXUkq27UjCuKNT5CKhDubh55gPU3Ejoph/gwtL1HPfVMetEPt2noK9aoy
s7HRLCtuFKpSXVgpc7V4whSIVdeoaVeHKrmnzYzbXzeP9t+HE9qkfQCrO+kVW9NaFReJCjUodrM9
hvFbHO+fcL/h0BmzlZtTcAuCeJYhtaqYyaMka8BNUnmCfzXmmFyoCOD4Rl0z0VeqtI7xkSD1kVqG
IbyUbA6aGZUKtxa8fvtwTSardCjFzHzqU94B+b4sZ/cj9DUQbQJ15OCySbdKqWVz3IUcrWjr3tKW
IXP2Kb9Ye/rLGUdZuQUfjnBQvSeVrWRChPqoJvpS2cSa3zATUChDWCw17Og39j8navhxGGRYqpVh
CdsuffAJC8bfH6oMR13qxYmq/rAACPRQMdvOzpbf8i1LehaEzLRTgbjvb+mYb9U7whEd10vGNa2G
Jde+J9kPb1nAwM8OZeMjv2JAPh+R3buJT2ghpqQhFnYd8rwycJXEzwL00ZXkpnMufvFLLinw2N+n
rLTfNvYZ1Nbif/1SAZwDAwPZyVOYbKqWNe4cF4ApQWtg4W7gNRCakkC3TUFFNmFRYpJmC8t8FQAP
fXhqMqLNoxUDIesyCo3sTRZYoEKYT1WX6K7BTUM1GzaA+ki4HCmC2ZpyLw4DHJEFlsYPV+LT88CB
PYxmjml2VpshpQkqPuOuAqh6lwOWjtAtr6Bg2oJ+j4Vws351oNtIl3SNO1ERQ2S5xsJLAHNXzGEn
I0quy1AbMCGkZcIA7PrLVgIHpULRhR9a+1mUJKGu0CrZxja9YZ7jCmHClLgHe+9LYpRBnvG5YC/G
6hw0qb2VPOf3EgH6xYzaLNFMiRanNUtGzAnAs4GNPNKr8kBx4ysWOylYYQP+ILZdwnFjwvnnJ5hs
cTtx4dD6wHCoudP7yLJSzsGGTAtDclrcZnITY0YJKu+mdhsnMlCUInxloZZni2XxAd7bKhNyA50e
hcYv3lWQVFJUtqCwHpaCWi2OZ7b4SrJNa6tmETQPFspg6cHp24k5VFESFLiI0Wc7h8k+cVGHyWya
lZ6sGZnr7Bgsw9R1vWkE7X6v2FzI9CdzY9E26C+qizgwhG++WfDRu9iuqA/IGXrjQPc2iiLpZ/jC
0HVzUQ7c7mEZBGQQ7NVYvQtr0/p44pxpN+YbzQmtKcCCHSVvuKt0V65y8ifFfyZQ+wHNlGNAA/PO
gcFmosnAcawJ/FiXZ4V7bMk6RD6kQWrYSSYYASdNZ2GlZC1zdCIgTxptAsVIPEqBGfnnXqJ9Jgu8
NJMuin1ZXcG3LLb55xsUTW1QQlmXxaJZze/vvKzu6w0brB4fkkwjrtNPL9HNPS778FvqhK/4qO3R
GXi8+b7uI4PXpdKWT8fJzaeEeyMWY0SdVnJYC09jAfT/Pu+/3CSTXH4r8+i1pCpiOVgNecoIz+Xn
Kj74qViCaVxKSLiVEnZ/isajR9BrKM8mz7xA7qQgqG80WMuut+o9yXTUh5oylBhpj5n9Isnd7xjQ
8Vi6JZNGDJSXzF56qYp3IwQP57pV0fFLxWxyrnWvXEpWDnMUTTy4txdtbBGiWQt+kvgQHbrJtmpF
jZCW02pCRO/vff30TSYARGhXPZr26QA8VOeFEhlqmpTz31CgPPYxV0bu3w0Wq1NgCviBlWpLYf9L
9cKiJroe51863Pt/Ydwx4ooE5eO/1UV0tNsr7UFR+B4Z4kQ3GNQPOhIH5WCb/+0qZ55yxOtEEWv6
vN9MyetA6HjgOZGcN5lwA1IVMXWvssQjMILkEQtePn45+MF2MSsiWADJ4CHjugp87UHK9H4BSWQB
+H3OYTrqhCl34i8mGeZTqHHwYtYFSTTkAMuCPLjXHz3d1QX1Z8ASABHlhbo6zrZnXkkmZ4fLx5Oi
bUnpqe15D6fw6xQ3N0k0opxQfE4hZ4+xO/Yz0YmE5Gbotbys2AoKrpwoWANrJska2YNTpRnWWmVD
EDw/SCTmZfW4O2wivmVyXjmh/C6GkxATCqz+M8XvilegWdkMp5L5BXe1GOG+1z5yNxtr+c+IuLLr
0ltpEW1j7EesxcSo2X5QQhsB8e6CqlcOXKV64gc5kmPO9/8vPRZhQ+V370lo47BO0e2knXztgO7u
lU7SbFX9xCey62LGvbFqAyPsTLY4VZTbvYgKCmMkrqc4G+cGwD7Vg2X55TAhqVkJnTIcWncvvtBr
jqsBRFSqlY1U3HnEFp1xtyybUdia1hQ3PiSY3pXiBUNRX/Yb9qUzq4yrht/WUKx21boXWVtFpmLl
nbtxZNYWBECZnrIvVxLhrdTDs7xSvddiRzBTPFNSISGSfVfD1X43KBS/NZU9ocLa5KczRW2kdidG
V8ABVOunFbt5yhOUADqLlr8PyjkAxQ7id484WRwrKamTNrNqfuTXZLAG4zSdejCLKmcTGqXF5a04
EBJmV/kh6QQ0ECTPQ4CgHDCAkbGldsxQYgDQ36AOgiHlUgwaAMGqknn0+gR7YBUQ0PVZ0GgZbMlB
ctXP4Ub/hzovTwnF3BS+pOWHSMcTkQruDHT6p+0p+qxyERAWo/iuMoy5/6bjjE5DipIrOgIJwH3l
0uQitfrL0IdcICY9IIfX+NgV9zJXk54FjpeRhp1ofi07KsvgkUA1LDCOLnS3ulkqfyDMxjcFwoLY
rVdP2bPeoI3HioBbH7MlBs7/ckfCjB2WQ2qgW5DTMBLsUcD6wY/dhV3rNvlCGwuAmd0PGpI86047
7AZ1zWDEQTLWyTssCg/ybZ1NPafeweoafSAFK011a3nyLCLQURe3CzipjX7yfaFJAkq0D+/NRQ+X
zILMgZFIo84e7ey1mLRUf6Sq+4CSzki6vMKxmX1P6GFXSju98pafTay4yvJbpHPzi6iG68PuBalA
myHdqz4n2JxrmjpiDsh6oKxb5XBla9Yk228EpQiRRdkzWACsB7H1fA148BIxJgkxyQCd+tfREBoK
17U7fU0Vs7JLFTOd5n5NKAGeM1iAJVDmo0D8O6bDun8TQnrHAyH5RFf3X+ZZTJuWFtEB1MyU0K83
tltL4p0XJYUI9uC4KGDUK+JxG4p6Iy7BU7LPeWul8gdNixwox8K9iiHJDeYBj1n07SWkb516nH8v
WJrdQgFWSY9rj1V7tKkpQQPdenrr504KmTykUieOptg0LLnpZx67S40UIaZhyQEFnFuR46+X+k9C
QP6DgPo05bRyp5nlD2YoeiTImnAlf0Sxx8kBtYADn53i/tTDCxIVPdj2Sj+w7mv6/08sllvFH1XA
4CvHbbL5qkH2qyzRVQm8Q4oFkLLFkfUzGqw9d1lwVQ5oqofTlWzNpTgbEENKYSV7M5GJD4pbjvhr
DWMiYxy8q85+upZ5rCtYC6V2t6DhJ0LHe4KRFSRLVO8i6Gis/V62nTBnjVvaJyZm/W5Pa+AZ7gAc
ttTT+qV0DRCcaCz5QY6TchrNT/KkZvQ+a3xdcOMNFx7Y2omNY4nwY88pscdPFhErumb4Vtnf0Ay1
PU1Mc9juOMRwC2wD02RXEVTscwvSq/FS7xpWoc41TXtAmmqVdyrANabK7BQBNj2tDl+4FZngCo5I
MPwdmlM39JHRYxTWsS+UzhAs41Ry/U0Dup0kfNknxsrmsAf2BXiZZ+jyL4UtYBShn+8iykkV/XG2
eu00bBzQo4bF1HcTyHFBaAGK1C5D7wQyk4Mtw70NbYFgcY8IwJNHNQdR2ksko/kQpt0nRbhTpEi7
gYMeRgpaF/pSuCM7qovHZW0THYQWTJLhrWlsRskftVhQGG07UMy0K50dgWNOs9UBzoXs7R8oGS5b
L89oh8lCv8RStuVti48wJlk8PqrbGU2KQd2h3v5Dmsm1j8Gg4wollhofQjJ8s7rMpwLD7NmztXZc
uOoHoiFtUK7YVC1YkPIN8yM0UnVq50pAr060dxV94lLE8+OF7881AUBsKhkUbt1OEZFKKPzi9ngN
A+HVGSrVtfXnC0ArXbKJNKGQRR/hHyVk5VjcT54Pf+XbxRJ441g8McbWGAVW4ME3Oxb1us0g5K//
+a/puIOqWBj9p/F0YHqZiRgXt6ldU8QLbicq+u8FVd54Eners+Ehh11d6l72vzAFZwOkryewECMM
kswuoYaArXf1spuNlNvYPu275GTA+5b9sZRAUwujiYoLlfBn8P3fhOAR7CavINwEwfS1dW640yrR
56iPfIKFcbitj0Ne9LFTDXNSVBvSHjgNWyU6e9eznTSNm4qPapTbUGVtxjVV+VABknzS8tWV6A/x
nyBP/6zYWdxcv3Z+na8O7dvse9nVtI4v35/qsYCuWT3Kr9/ljLtDt1U0MHmixli5UK0FhkF75KQo
MQYPw7KVa0hwUzQOJUCzQHgGRsWa4CoqaicYUvVx7eu/ExRdREP2NepPQUXUcpGmoiq8kmr4JyY6
k4F89CwwJcdRxMrNg7z2L96gl7TcQszK/BDhqIGSTK8gkzV7+gKPCiILKtuPBlJ25Wk1tMSOYrpQ
Q/8vO3ZXH8ogR6hyf3bPZPsHy8d0WKSKTcr5RM4XVlmKfr9aYm8SZeUpKX+9nLAxdLjF0tu+OkSk
b+WD8P0irW3hDyBwTeC+XRYjfp21W42qS5eUovgxEuW4Ip4HgnNAyTwQwkItkZOEltjs7O2eEIN5
yRWVkAOQQ9Nxj8NJ4+pu0grqpwKEHeX44sglhdnq6xVXk/wYRY7M/DF+kZIwWRayXbHmL8ZteyMT
QQfsh3D2X9mqJdqgovjKdbNy91yO6xLB8btbkiff7Rwfa9oVZhHBA6zsKAK1vbrjXg7GLaioGzCK
CI3qEezOHfMSl0jRFCmMbhizyWGLDrau0ZOj7MKf2EmPt9pl5BrwHwDhvRoDYouQpyCAhjBKpL6j
9vSCS4X5GlrODJPgeBpIurO1vfFiC9Qst0+pKM3mOd7MuONiRIWMQglySjc3YXIsmYtscZ9o2XhH
z49htULoHU72Uqh7Qu0m+UCTJkxiwKqfpghBikJODeDHZt+MzMyCWJKZL5hnbCPyd/CUbUuCzn9V
O3UCtrNx982XIbljgiVHRPScRLdqjQngmf1xK+/TU+0H6DtY1k775KVQM/z3lNi82ufI2vQ0SV9K
GTQ5bTAp4XUSTaibcXJPIa16gLdB5AgJl9h2JQvoGN02fjeF7CHz2Zhxc54UhVIvbKkNzkolPMNU
agbcl+BZN6DdAuKhQpqXCeR1H40WaHD5Cx7x+7G/HZgGrHXIoT4OTQSlfsNTDGvX2KNVLbfafRs6
u4eF1QCc+oOMLu3Bikt+yaE0+e7LDbwGjXBoqLmYyXvbWjPht/fRpFbCTrpq8RpBnKDjRsFU1bMF
zQsWtIiT3t/4jByUPsfOOWi7HtVsnpOc0+LVmlcE7bjQG1Uer9u/aDqzHop055MIL0m+5dPzUU7S
t4ttg+38KhEmnqqE0E7dpu1+O7To6SO6VtFBxM/yUzXIJxqJ5qiJTNzQmEX36m7MXGHtqcCH3FAU
TUke/6cd55vbEdMLV5vXS76NWYZZ57Pp3E4RCusiUepNfPsTG8vyoE2TPoHh1Fv/2XOB+qNxxmsq
LOdzLWaFqWVq2OItjvOb/QKlqhG5AwizqZoi+Zy2I1c8teQJzCT5d8LsSg5cBOCnuHEEZn1kNUXP
u5mYsUmt0PGBxno11zM5QQQOEmodUDbhYDk46dTXUTAJG1I+0u9bQmTrUS2wVZ7HBnL/o7LbV+Q6
W8bCybtMmRBbp/R7JAD8DvxnGBtqtkhsBVFoYqKOpCjR5WUdSrMX6p8/H7WkANXKvRmrjTV41kso
mmlSEE7Y5WmrNOfUGuNce1nU5Xgxx8Yb8r4nn+sqnWjVMATO+p20pTVrSabutyAqOsl/YfkqXWMC
xFL3jy498SDq95shGAOhDuuXxPxxW9bNNdmxPLBboiT1yppMF6mLyqPLVskAFZowRQ9PGP18lKWm
eb1Q+AoBzpPtHavmdhuf3jHQfzgL2srljdpCyZ/ov7sXeLac6RaY7Wyg+SEnUJZoc31wf4Ctcwwq
CcQtQrDrO8UOg0A2pUVgohEOopsJXR5hhMz9rSD3twepSl6cap2zQ92XcsA5MbFU3IrhjwtiuURE
1OB9rEJTwDHPzx0stbHR6L6XOCmNOv9kSDTK+EhNmwAfv4NXiqje87wcE0TIjMTBqIQmMYucFr9M
a6Q6kaGpg0IPfk72gHS3h9PZZ/rQxvGmj7PhAdHcvkGk8xgjm+eSgz5mZc6sJn4idjMkmpLyKApn
cMeHwEKCgUXSpZX4Aklm0FGZaxgU3it+44gI6m6UMPQhitcuvheMRtxrc1Fxmro7Z6lWW5Km6TBK
NJ/RUW+rCwBdapW30qUPDzNYgDDL0t5ERU8hiiBO2VlFHAc3yHkYYdTmpESRFt1t21+iTEXaBSiO
p+3Wi5CzmZzH5BWU55D9Ao5Jts0eaXGJ2xwFEaG11vor4N0O+GPhCmTX+uTh4eNnDFDYKgv8uEoQ
4lWBjrumkj0qESQTTe9E7vx1QXUJrstQtAMx7MzaWDFtaiTLMcoL6fAO7BOsrUPfzpc4+tBiJ50D
STuTEm3XIPtJ8Rfvjga/H69SWd1t44bQgX+5ruNLP0HobyQFNqSrIqMXnqhZH1sI8ektYsHB+FCt
mCv9vEdejMveBw3jZPvm2TMWV2S5EgOSU44aq+WO9tiZGECdqCyil3xUdDLj9elhP9HdNEMAjZOl
9qmdVk057gD4ocT91fHB84rwwEA2lQtEmKkDfwisiRWIf22SvhBJ6jVl9krqAmMyzCByCWXBHULh
iCmulAihocEkPnsIjD22QyYIQ+684V70Xy4VJd5HyFnmthlygpD+T142tfYG2X2ApwL92BZaxCDJ
Z8WjVyTIV50Ffi/nUjN23Mzc73UdB50pp5VyIDgSkDSBBVQGxsbcgavE00GSq2Ee8V69xY38lWC3
le8oEOGy3+qXWpN5RkhmRP0P9Gu+5TRaCVeTJvWnU3Y88I+aCvpJBW2ZclGyIt9EpnFiy2wolEkh
KWJiwNEfKzLkEmHom3vtTkjabQhEPZqtUbqOA2OJIAodV8oDTZwxlmz4AZY9DmpUO9ovs8BoaUGj
BUsDfkbcVuU+ct5lMU+WzTuuIgJhOQWiOFG/tN1gmLGoYbWto3VAULT+kI9fEo53iezWjJaFNhge
z9XZtiLu7UgNCseV0mZ3iXt/eQ9pQKWK1Mwl6u7HYlAHGZ7q8ik++chBs8t3pt00J8SN8Benden0
lmrYjkRLFH/x+8h/kSJnn7j9OsTGpd+e13+LqIWWistTWLmMX4D4FdXhVz8G98pX6YKROk2ASwgh
t3gpJLGwctHLGlsxqfv010CmG/QwdC+5/AqW4Cm8L0DsvMrXTecoQtjQ11WSQcKATVJ6TY5lazdk
HqJRLZoS/9O2LIQ2m7na2rlhDH5rsJOBqpU3u49BzTSptWfXqvsvZ7vZ2eJHZCfkOUxQnEkmyQAN
au6AmxLTCF4qy3LtqqLZBOKP81d5jweOlT+euw5ZNi8psHa/Lx6Fx8jqs/rPwtlpJBlqthzhEGd5
FAwDOyZmR8V29auEtD15ogh97p00UwSm8jsdpgyJlgkqGO4kRo8bFu5E0HNjxwcS/kLwZ3gOPkzL
YTCJk3XsjPvuGzA0c7N80YCsECksdWEX9AOKfqr6hBssSg1pXn6qQeDhRA9mg07nKepoa3irWtn8
lRrsmWDNUhtsiuKenKBusTc4W5kOXJNrY09vJnK2hVK+IFL1gp9+lgFi9y7MmuLDozmfugwnnXMz
gT1+JsWscZG+rpXcGmtCMZQ/o7VM3D/Zo/OPkiFEOuEUBnOBxMb1R2FbzWLDipYhXezfkSxPywEI
HC+ltmr3lWWc06uuazoevMlMc2k8MrN2+fWAH/H07Pv0UEugU+KPRZHNe0FnL3sZ/vr7H+WlqRm6
GR66nAQNg22ilJQmuiQhHflQa794cVzXBkQK9A3T/IMQl0tyIKihkVsEBhzUWmimMChIv4IhCDco
cgjrzgo2Lst7AjvPZq6mE7ERhJdQp8FzmjXqDCjxx+MZQa7ZD7ScOqj1jFhv8LMxltSNsyHrSPzH
XJclCamW6qyKdiql3EGY3HmrRo/P/PQYrRcBXSgWqKtLyDZzIiBxOt986qDckwjV7AuovGoBnP8O
ljSlWr50IdruAd4P/fsa0/LUv8X5o0CiulZjwSRnT6rdKcnx5CLfH+noCS+ktz28qqRHPCsGfC+g
lo0lkZyHKihTr70Zumuve008NPwSlT5gT+ta4yHXVSu97eRGV/jn4BcWG+cc8XFvVXM9q9j75sbE
iMX4LkE+LjizpUg7I1UUevHTQBi6++xo4n1y567Y1GLbXPT2KIaFbxMWF9qmdGrunPUYoSiXAFih
Bzk7MQKBXx47tE3p/0zr7WlIwFNcontvFq6iQNN3Wdb2JSf8kseAyD+Yk8m56R1FPr/F1+TB0bLA
G7mh8MKJioohCZtmJm/winKWdKVzPTTVdZNCNVasGolWilMuzAlD0mnmQfdHFSWGGVy+XNvfZPS2
9W4/8JUz6YFukmRi7iKh4VagwLuhrSl6tlt3f5GHL3pY2hZMPwVFFPGHXjs78GXAAqA268fl9s8h
b9bI8ZeKdyuf8MA7OTJJQhAMaMVt/72djAy/z1pgROvbYa5Op5jdBrkMy5fwQajz9lGW6N9ItDCV
3LhQCzQ0zWaw//dz4sMzZC9PUEC86eiSk+Ljf8m4uLxuiDGCubXaWM/jDLU/GkRjFerUadf6fSx6
meAjuZncBGnb13rilN/syjpshW38+oIroPEA2WqF3YRfnKGTJqe8F2pP76b2HaByNqlfR718vfOb
Ph2EokXQjsSGLEdzfa30UzWKq7aLgRKMXN9Dzl4GMLf/AELdfS3+6acCzhO6KaocldePlZslO+6s
6jfo01nwa0YydOTxVqreI3BudcD6O+VRY9RDe3m/t0ZeVN1FdW+LIhe3LsZhY69ysDsGK6/PgVSq
Q4iBiLwbOTfd/FGYR580MBT6vsu+qBSUGijvGzlzCh24IIEfnP8BMM8IkWvJk9OdzMuPDmYJ7V/M
WHSUvCHKcc2XudG+hZ5j72VQoGLynwWlgIjnNXmVoiWleuVuW+GmnF1874lBPLRVc8JIhv1mXJbJ
ubHli6/Xn/HpI2G7S25PeK3KVS6Gqi9T9Hn6kZYSVAzF1lqwL40EmbBgrdniih/15e0sp06szgPf
wfdkpEnvEXzoDFfjUQ0t4PFLVg8UCXNWW9KSQb7R7z6Q6yMxXyr3IKinM5g4X2ytrrLhs0zh4ZW4
xfTsnoKxjvYmNf6T7ZquVGBiNNselJ156NhAguZwVIYnjF55+/4hCsj9X6DpZ1r6WKwcAivVEilt
iRRWKtEuiCp3L1HNb90R2Azo05kZOK5WBrcgskwXnbBhhBN0+mTanyQSJV72s6Iegw81u3U8bfQe
ilO4viRezBxFIXn5oL9YGtdYi/SZCHjxmOdkpJcWfOJIvVELGX/RgtNbgAvGeym8z9cHfsRXzmgO
b0ZP1gvQh1MuIb8/14BEz2tIcwiUC1y75JaS600sLe8kxi85pmYWs8d0TiJbUniNpRO98Au8MC9p
aqdS7df/yianX7fI8Xm2c8wi05oIbic4MGkv0J00aVwyE4Sb+uaGyZlA5b11UY75kFqYpL8+7JHb
dae4G5+yw/BAS+sodbxYNNrfhtdN/yw0EW22o80vTKdtvOe5gRBlONVlDAS1bTNqaf/uPD0zKjEJ
c73BLSjLomSVCl71jijVy3o/F92I+lO4K8bwd4vIJ3/q840A8Dr6YzsU1ffJqwHiQZQPJRH83BgI
13VB4dFfXOdYmfFpBX60EdF9Ijj8uYy9l94gIjQNSFSKliZDyD53GdSy9PUrt3WJoyspP41Ce8TG
JEjl/ShobuDq8HqE4hqO0Rlya8PVjNrq4V3QTcXFxI34k8a+vv9DMQcY6YfU1bMaLscjZ9UlPRBf
dpMJX2Mj/zfgLFmIsWsBawLcM2Ivjz46pkeuKGVY8fA3HuN53RTP0TLB8ly3i+fdPujKQN2z8EXq
MKohecXoDWYM6Cjxs5uG+xmJilRnjfHiDVq4ieLvGIrTz5B2i0go6tnmAfyZXD6hEu7ZC2qSiSFJ
7kuEiFJqbtuA3xMb3DmeDXtGC8BzyAgb5qUNg5kni/xCcKOxFS4ADC+u7f3YTzMyfflskkOhKtLg
8NYRDItz8GDHZIxupJR/hSJLJWi0WN3oIfIVTfcojeQPe2+BIxsXbdy456PZEhOg+rJe2y4FPmxi
p9moS/6zRvlrZTatOjh41MWVXq3pjdSf33eS3JCszkaymypn0yGHcguRJaS9Jwmb45s7KkOw07eV
2exC78ISDobGWtahyTr8om03vWbNXQzwHryZ8ypcsMxZfK+yHkyPeltgePS4OYkAxmk34+l4lqLv
l29sQDc0R7nfDP5KCRfqzkNjVoBRiI1+KIDOXkoAFLvuof1JfgFfnHk2BuCzFoNPAFXwcxrs/1cI
T0J/enb062zLBfvhcH3AxYtRa4DQ6//I+PWlSRBuBD/B6JtCBXdyYkrhBti9FTouYwoBvKgHjyBk
28U3qERi5PEX195TeohmycurJWWzDefN5CHLL64sw/pwBjP95xSeVkEv7Y7tBW1gQYls2nm/mTMU
7h1VdLJs1lkkUecJMV3L26IggP1nN89eljAJcE1P7Vf35A3eoUAfobAFy19HdRbKLXegPCt4mBM2
wbcyjxQLYkaNfF3F5EzPJxmkFQIhcfvJGxOio3vuKcRdeyxPHKz1XRx/NZkL4Psle/WcHJwI4E9X
TJ3tCu6nhGaeTovJo2btRVxj4o2P6V1Yp0HqTo8em67sQZkrQJcI8vmhVdb/pH1ifcA513fCyGJy
aMhw73NCqivCLkLMPJUHWOsVB8EzjDYLEW8rhIQwzGc44HyQzGaZjtVXKUuQF/58jSTmV5QIjyfE
2nnKO+raJvc40cmzcQ/GpODyIMgcxWfNyhE+yNW8SBnXACtr/EaihE8ntWOMIZRs3hDtzFGyEYlj
/Am/RAbj7Z4JMvciOJnvf4UZSVUXm2vQVpHQcRE8PIMGr7Vgyb7wpKKF7aAJQRNzBtZdYety3IMj
BcNyUAmPWGe2UK+LatZ3WRt8KUqp7PiN17TRPJzeLR7Z/0q6bb5QbpjIeXsUhYqfWnoLSYRTfP3X
sbfyWDjmZj3Euz7JyA0jxKV8kbgNaYESimmFX57oq4cH0/6OWq3RRGdKP2zn5x0DOf8qUKKHV5/P
7/k5MP6km0xmEGEb7ufkNFDVJ25B37SHjGlfkofftmAUn9yFuXjBM3GU8OMzsgXbHBwVTq/SeeS6
4okhM4AzS1w9TiB3LwKkBCcMr4mSy28W+yHuRXZnNkjOWl0z71pLomImCZ3HpcUqgObzCdQmT6Oc
/7WBK+7xiMOcrXu8lGi5Bc+2ALpElnF+8+PrOqiv3OK7Ozzg+fo5Ix8RKYgxSzt9p4qFFY37v5HO
NM3XinumfgXoC3U/PjJUs5PjRDhlTjPwEt4Bljdxhgz5hm+FX9aGfLlagpVoz6xl/eTMBnuk/XFV
YKkjlMdqg1WwoEVVG7zecbQ01i97ByceqCnqGQoMUPG26cA5IO0K73w4XDu9FbLHH5qV2IExZBmW
eBavadIADElCFRgg4Dh4EAwIQFxO9wDBruWrUKCOGeAJ92EMEZtivxoiqcgM90VEVzqpHd/aZEwT
EDV1BmJVzkUl6QpKvgMs37Mxa7Z1E+AgNURPlQa2K7TMQb3d4TLXWD0wN9Fmy9HHPWoy3JUTlmPO
wq4LdhEVaPl5IVJrodjlSvdzZ37jkRw1YDJ515rr4EcxLL54JKOMWI2QtJVN0M6peTa0msS6NHxI
xXb5gghbyS2dveq7urmFIGA8761h60P9qHlskLKL2jJAsQ3mV2cKJMYlybBqQrp5RVdqGU4+mgSO
HPS+hogWtqHy28t3Tg/mHRYaHKFYur7SoRDnBUxbIUcyVRIaTtxYT1t3VZFKWJXqyCMPlCTqFFjw
9tiALCWvauD+jnq0vrL4btcBMvzXEH375j3jjx5WlUG/VadjxAvmulcLrpe8ns9yrzbQ40bwIM19
npq3FSUjibtzzI8vfsziXOjIu0SNIHazfB81w8vTe0cJpD7QTbPC//ijeM+jJNMRB400Aaa5c+dT
xnif0pHLPW2HhZcdATaQs/ZGnAgftcXAeu8xlu7eikzQSMhHGnJqylN+l4mCqhPhRRTWvrgmowtu
FkIP5ypi8Jy1++4KAJWL4wXf7Nbf0pILn19i+mGtlt/osz3p0Cv9Urov2g2+3dC5Pi0VoDJqrxXb
Z5NGLnj604TC7HMZdl7oD2b0O+JZ82r3iqMxWRSgr+LXQg/yokv8O0Fvi0g3I6zOk1T8UsKpaYPC
jfAvfBmMn9Gi7e+0WAK3NR/v6Pg1Ig3sik+VddTZUO/2b/EEiJQPNbFyVdUwnJmIajSLEhxPsRTb
nX49hVTqbq26sOretZsUi7WSbvq4XAfqeD2jareBi/0FcXOWhLYLJHeVwC/adkvuozTQPyLtyOPI
Js3V+1QJ4H6NOxApRaAj8w9je9kKCY8HQZ4Ifu3pghOf5xVLRcIOfvRgg8vJEJtVjqxI825HLgPw
IlulLpELO0sLifszfUeFj/t7RwkAvpux9S3Ccxc1Wl8VOHvidgWtH1m1A1Qvp4JUjK6wcqK8wjqz
ck/7GTEQBYZyWv6ssOWcjqZYntv1k/174/kYn+Pi9UP5pxdxzA3NF4RfTNiAsOZvswJWDXIel42P
c99NrYhNI9AFe/9x2EvOaCu0koTxcpCAho1FuYkoLGeEb07YojOHfMCUIL3T83M14JGc/GgOY4DC
soGkGJQXynukHQBGS3VKd02UhYrtpYrDe73NX9KZkae3+n61v/zBMAgc4WYxOYHlZzM6sfHC1Ez9
XovZi9ItZBChk00NTgyG9QN0bJmMgjyKTxmVIjPzi8QKqnda1xDoMpiOxpIaQBJ61KjttBjDg1ju
dZM/Wt+5kj38X2L2geM8pzPBKGorrSvIN0XGRkYdRKy/jVJiYaQa1S6oxBXEKloPxwnQgtW8pc22
+rAZ3hPGZ1uTWcpbIvLto6BiFNnVU5OF70el1jzi8hBOmWrTu6eVxUIVhmD2aHcsiG9r2ZbGS9a5
VVKYHe7BkjrStnqdggrjtep9AHt5Dns/cQkcdvTeWmf/W7jSrDImdlwueteb51n5Med7qM+9KuK/
4EhZvUPQxJN7ufyBjkiBDwS4u9nxFWyD4ckKPW3kKgWxGh1966RfG4zCHu8GdCvbfVRGrNdPdQLM
SKscDVJMz9K6lXmMWJIvUyQWDaMgf4mU6EB9433YarrVM+XrbLK+gjRNac23pR6s70QLNcdloTBE
EcddwE8cI9jl67rSsFCGEB7x4Z9mIER9FDvqc78z2sSzQSPQhX8w4jlKNxvVGIBjxrEYx+vu+dYH
a+hix8NzGJlx+gzbo81pDjoc0rvQtLzApx9qugwxO/wWe28tdnP0zuLFV9BNjrBdYKCCPBoaZX4l
jGArukEUvZYgq/x05g/Bo/cMlWM03dp/daztjAC4JgN4i/4GDkiSd2I2IYFfWH7kJ+gEbnAYTAJC
QIwITV4eNl1QKtSya4JueeSNuZzc4tpHYHAukjjNxAVUw+p0f4wOBbBVgkRnA7aMFecjQ9rIrMrK
RW3LIb5AAQLCnKAIvc56H+Ze6TPTjq0x9nXM6F6U6WpYZSRNKStqZBwVOw5xX057SlSXHnsQyAtE
Bxc4OVDlYfQ0rSC5IbgrvncG26dj+4fGjMWb3TWt0ktz8yywDTgVBjgChyoA7Y8XrMsszG1Dy8ny
4J80kNufvHo47Hd1mkjUKk74Rz+1pg64t1ubF5iUgqs7W1nUChHeHzolJLAkYYj5UD0NUIO+Ozmp
G3J1HCbLPJlNevMJnmF1Jlpa/RK/IM30sdrpthUVpAVcwPmnwzQNE5iVDGVgeSEo1W5a5OHsnn4q
9MfRC2Sy92v9pQ9WGtZJI6vDqLjXnS3zy1Jlyeo1fuZ2sGbkMFjCrNTt6t125TZABX5xIlShAFwr
xlAACA8YFp2tOIRjhgh1f4C9Ieq91bDDHG0/83hg1Rob/ZzwQYzqqHelya+l7XbZ0nRHhi4Sv2KA
VP97Mm9JGIxFHYfDQjJq4PvNVAGf6yVTE7Ph+FHIzoxHKgh8RZNE16C13pze5tpVgoaPjh5JlBwy
9r933jWoPKoPYVCroZpoXUu9w1emdoLByBCpSJfZsIP+IdttFnqpbSP1QLuquXabBLT9wabpgOQP
xeXkOs1Po5vN2bD/VR42uAc+r9zeVSMKr55CHKrmk0rbEQODeJX9qbDCwFSYRl9ScnotNIekZwNn
HEOadP1oJ3ZTpgNrmkGpsHvClaRbRbN7AbLShChLCjWTVPY2+vEgIfv65KPv539OleB13u95yIt/
nsWBKPg+MhkP5joxXWQTZm+mrRXbbOa8mEmAa7sSAkPEn94mXrN5BGSWiGUqOsACnpBTa5bYdd6a
yPB/pZb/SHhvz1zgQFcsYFiH3ZBqcCyNjJ7nJuPZarEqZcz1MHsWIEu38UT9zECs/wPoTNsdTRD2
PI6W6sP7h5uLOAcl8cfzCLCMxRNOMq1EXeZkFMnhoM6dXIuKcyG+kIF9ZGNfqpaSNk7Ybx5JTEV9
mkJ9iHbxltPnUjh5xegp76+sShAUF6nVSoFbB2HlcfIuJTRXhbX40El+egM8bhMSFSuxl2Ralhby
7XdnJCGGHFFgOSGdl5PxwWEzsRtyAnocUlMxBdCfmAxjnP2oizqpIB+d6m4NQi5mReUZi5dGWikC
E/y1ICcerE7y4URyiOjuWJ65omm9USU693C0sgggFdiiLzijSevgxI1N0hzd3gI1mkUjyf8i1WCe
4vt/HKmotVpV9r30Yhh8aJMT8WDjizHcUzFWxWoUhtn92NjRDnBkKydG7qp7z5/xiFw5IOy8353r
PTA98G+t4wX+ra74C6+m7KXoVIdkNQI8hnwbrVMMbxKfB2kY0/S0Zyp0U/bYWCssxp878kn1salY
KmC+bG1ONkxpyQ3hTtHDRhMTgIRhjOpuO2mOBKL9RfSKMsC5+fIxVilLRiWC5xK5uulrvgwWmZgq
NVJoYyfsVlEMu2Jg1kt+SwDQqQ4fnHN9EZCATmjKoaC7fXUg1Of9UR9qWlDbPUDKJEYN0Ce4Q8D2
bkH34rH7+OgoCtHIXe2UpzyaOy4nwoEHLu80wHuU8POBk6usbPzLHnBAJ6Fz+L6UUWGayafYn+Ze
j0eApTSvevQKlvJlCSh0popE895wO5JMS4sTUIV5NXc4krdbXk2vKiZ+/nv2gJtY8T87YIkMX3Cu
q1UetxKRLIaIEmyq7giywSdrh04S558n604d6N3vNpf0zUCcP3EXNDJqNmG+ClhmxkhFqbi8xNC3
2tBkzhAjPzNzIhZPCUa/pukgnYD7mlUobickPAP3FQGpVC9cLTypuvpSO2/vkG8G0eWIyzg+ClVW
3qhVL9acJPlcoxyPIt6G4pluiw9Jly01y97H/NXCXG/xkfEomoysrrXHXhqsvYOAwUJzoyO7cyxr
mI6IiKhAy0TUmw7y1pDSC6OJuIjTjUEtGcGrldQLA6JxAkxm5fmqb/hFMrHBKGFfsHCTMCAvpBF1
P7+ToD15RDlBz+PtqI2mVP0SkdUi1Lm4Q1623aqL/ZXa8oAG6otz4Zdl3yPwYK0khqT5XipHKje2
4gTlRGqBqJEn+IWpLm1eiAS6UaVzyY3UYTdgzUqscamnsTgw4T7CHxvfzKxGjt688ZK+qrGH7MWR
doe4gymdL2UX2F+pCyw7I8KXg0JdACKuUaiNjCnmjZ4yYBL30KkR9dmoquRHFv8sUZ5zuFyprvCn
NFDRiQ3AuQJlIVIWaiD+YhjQMd7oi4W8AUICJtzy6Lfsn4bvkpdGAzl1IjGGG86xrfDvNycqCmF8
lqcmj5EtNZHM/UJgnuufcdSF164UCxDMumhFKPDgahlLFeDBlkbVyTwYQkmuFU0UTAILyxkr5vEQ
y58fVpKgESfpZ1d0ey7B4zJwhPWi9BEmFaBB8Nz1r5LBj+uvZHcPwiaRre2Ck48YpHnzZUfCvOos
XkKuntlqe21pRBo2iayinznTNJ0sZU2OG4NCD/fB40gDHon+S1mP7bZ5KqEW8Dz03uxHwe46Pp11
GFsbC8Q3Fy9hhls2u4ix5dQbd0JCKzNBNpzf0aumGtcfvQ4e8Vu1YNupQ3aYlUBPErX3wmG4vtw3
sSTnnj3xcK8ZdVxwHEyU27pPer9KFv2HQ/3OqO7kTelqA6t+ExHi6PqIJvVYZASllEWuxOojEDe4
f7CRefj3UOI+ICz0NkhpSoxc7yulfygRF/QXZJxgOEmaNAPFQ8rm1sNEAV6pOaDaYHFehnCtgS6f
BOeuTtpgje/DPwUWo3fE0R4bZpbgT5ptbp9TA6nhxDX8PimdNDgdOf3ZKenXwlngaqftZl877FsB
EXIJaFrK/2VwkGfiRWdl28UjDdmv2yJk8PDHVZIgJ+5CIGaU9acN/hkGODy5wKRj4XPES8c3WT/5
mG/cHb1ArSQJax/pbIMAO+koo1H/fHa9uDJtpQO3bcgSkFTYIEIEcAX+CRPMi5NHEjOXAdxHIwzO
UfHpMkivrhWIL/HNsEGxoe17jLA5tQ+Apb3gRYmFQQnesYxMIXBqC+hF7wwVrx4IfwsDnqqvIQ0i
eBmoUX3JHShVd5XAx5Zxud2KXwCfbHeewXDVrBi3F+msMADIfkAqsYr0ERKTv9FjgYK453kiKc3v
OloSXQpllOhJn6PTpFuR1kSSypUvFa3Se1pvVcZEMQ/BpvpiIzC8CbLOjDJz8q2jyMh0KphCjdZp
JueKjhhaPOm91xSSXzrsp6WzFQb9zDTonFbY+IIfuZXxIXJJ2O2gIF4yCFyWm8uPHKd8ucMhIESe
NGBxKe1TPXUONWMF4LJ/kHyfccjFT7AXSBHI8unUR1LpGoHvf8ns45Y4LmKK+jwEO9tneYL8GeV5
P60b2+XiLR9AC0aMT04opnQxuhQWEIq8EHs75UYTard1BJdM9benU2i+hNPTjzHcScJs+mgmC66B
lBWOz8oKkPGWkgmumiBD7s+wOT6Up956GCKNY14r+1So4Gg1OpA/lY6F3gbdhuvBuaGSGXQXKTos
NG6g9bouZ9LUBThcrZcb36xByO6UibB5HwuvJ/M/40qKxonh0PAHpXc6e3SBdHf60UcEfiD2AMeG
7qxxKa+N0wLl93LAadMQ+sZn6tK+0i30CUHFuDVU1v2oJhYlvt/wxkivTEgrHP3E9D3a3ENvV3Mg
SErp9/5993BI/OzSzVhDDH1f5uzTqpA6jmpmQKVx0nO5AA/EC29BuGYpIXvgRMxPhK5l/tJWy/Bg
nk6hk2yCE2gsjKxqDALRAdyMNvmPBt4TcahFbsTb+tcC4bIYQCv21q3x5FNVqn7GvEIb0f/htA6l
MsqDw3e/k1I6o3xKWqD/ipJqEnhuMc3ZuAhpeqdmO+Js9BiSoVs8nsDcL1Fs8cwVqrQOGH3x30Fc
/9hIeeHhuHY5h2cZv0+R1W5oe6thoW2yerWEuqbKIoeCr5xKEKxFFgklZQ9csvNjPr9LFa8SWbHV
iDLJqN+0FcXad7QXoe4mC68ryjlQeoWsPUnoBUGKe0ou8IGr9QgkONzRnlBMpNMTeorcDM41TQut
1uTKseLspQGrQNiyLn8E2SohuvgkqUustoGyl+0WYV1fTgfi0GbBoqnUD8jog8OEpJ4cpAqOHtGM
idA93Bui1DYExCP6P8j4WuJu9TPrYKFSmYITpLOOSEopO2UTAxMb9Oh4l73MkwT7OSi2po0KWwcH
iouOe8sxCZ8rlXl7qI1FEpGBA2d+zTe6z5TPG2VzBzjsSqSgXLvMxk6j+oGTraN4Xmzkv6QixUw5
CwFuei2fW1/1Dn7o+RyJSIChrzEhD4ybVCXlt6NipxUiUZPLays+tkOSPVeGHVKs/ijeFJvJLMPm
sLsYo+4bNrc5VnmcpAER0rdiTQyQHjrohMYiqEBTCEBAKcoWXSP+qG1HerlC1DMM2qhaPcj24rtn
MThswA9MdtpwH5yO357LpjHTIKdMe0MfmBBFyD3ER7lZWig7rmylp1wIygsdje6g6vWthNDjZt0B
ADNHRSXioVeMgN3LpidHpakapZlleN8sXvt3aswAexlS2UzVGWUMWB+suloSpzP4lZvneGx9FGPR
vH9l4iDKAf/dtgK49Cs0r6EhApySEu0yt+0QPmmXFx5LgQ0d3DmM2GtgLkAG6kxqyJveywq/gUz+
V+0Ubv+xHd4tR19GZRIPnVyOrnd85ghF60rjGHaWGmKUH7pDxTFIJR5Vmox6LqjPSPRNeC2Xftj1
OjIbY7uWIxEAg5+sVts6TVuZ39NV0p58gkqoq9AIHA3A3HrVzP1iGgDfUg4XbyN5tI/Zy+cQ5T4F
O9kLEYNxTM/fngWaaiAs9NQMxtSTuBs4ZCphZI3M0OL/E5amtQWjxlUxwGe/sv4jLZ3k9zcMNyAK
K5FxlIRv3ruvjOoN3nZoipkHnF3kDVlL+/QNZ+3bIHGqZsyPjIBbcY9KUSYc+aEf7nFx6ces3IfF
58w/Ju+495vhV6168oz35IlJU/gHZZN6hU06pOoJXhQp9LrPKqZEVQKpYal0VsSTWrBr4y5HXK44
ty6GHh9O0s9lXEjuk6mg0KkhX+QwZXOGADFh/H7jS/nPZEKlQdw1raqFhOLqVSzQNvjBLX2kUen8
LHnfCtbJOHx/WOrhlhfF+/r6F79rJEh9JI9YhC8n03PH4k/BPJ/G2EH5AtF3XZdJQsZt6AIttFY1
aP7kIbTPWHc4QytjIvAwEcPp8bxC/8Ya4WG5zcQsCSwpFH8TlpoOioIHgx+5CEsiSw68m+5TSefb
yMXj5oIZkyuhWi7JkCveYoK+zyPBXZbTlYEX1qARc9lZh9tHDdUtFInxGJqNZZhipOlFl5y/AQce
+T6a5I6zCOYeBMC8UgbsOkMOnG4sFT8g0GVUnwX8vC0QefrpKZMP6sxGMgTdYzWFnLsfIevcWc6M
Km68qgkQGt6xxQ5Qg4O8nWgB9RrKQSyGRjgQFGRLD+RRzUqojemOBq4vIDleMuKnUwmIWSQ/GyZf
N/nBStnayZIarMT18CVkneyYulL2k7jbds2F5bPh4otimHdpY2SmsQd534JLnQ1Rg14rjNk8UpiX
472AXMf2EkCRhRalqOu+lnRM3qP+81TmvlSbdtlf7lWemlRXMQgVsST5KMl2UeQ6pOw8/k7zuW3U
9ldpxi5+nhdlwFQIj1kYbGqYj8wkpyYfIl70EwHC4+QCjpKsSBygfmYk9i86SXk0KuK9xZ0+zUvh
+mf5bRkbSZ0e106qipKiymQ8iXVM0iQe6ZmRqaIaFjNMEQ3SfPzMZ2iZ4td4vYXxFxx0BsGgMRM1
pIKa3wvZGjZ92Oa8KQYxRKllpcujM7ewWpzjoZ+OsrieXSwadQCfGFGcgr+pZr22wv2gl6mGYk3T
sHs+jMXGzYR0ANITrvEn7h4nxcTY9yeL1Bqieb8XyI9fids6j+IlsnZm7zbL9ZgYpTNmpu09YGL2
14CamwKfpLcyaaZrku65vt4Du7T6Q1m/sAqyjOzjmercinyILt7kyct3y6rkxeflaGELq1YqmR+h
JO6UBZZjNeHyvg6UcuPzv4tLYGcL/URfE7Y8h75ONe6Sx+e2DzPdKxqa1mhJ1IPCN2kcruXclkv8
081oc72XsPxjfDnMyba5lu18hXHHqfWLHaegojJuUNKCAyK4S0xTKLpyVpQTWGj9O6LXftuQi/ca
U8+RAEBdZt6gTMziI2QG1nEh5VpKe11qGSRML6eIzfoUmkoPXqnRvEMKgFX33puCjRF5cGiT758i
QmG93BrPPnFNNFGI1/91Jd+fRkMT/7J+2YPDRk9eXFnIj7Czo3Omu5Thv5kow7NeazznZ+jPQ/Pf
waeuNRq8wnrwR2si26lagRCX2GonL6XJWZbDqfVSyRinLWyvKDzQuVnO11/er+YtS5mOTCR4pxWo
ThbNkrVifPgz8UwiyMqOBqSyJckvkw/cC/wde8OLg8GQYxGYWgcjzvoNHYs5a0sUGlLOSmXRYDT4
8R7BgvyzkV35bsCNgaAB2Etz7D3M4V1CoAez1TTOv55EkDPrU+q3BIx866lYk130TZBT82Y1wHSY
gXWv8TzjaN1n+p5hJYsl3GleVW2sT6Edr3vlEi5vNHUsq0n7v42nYjnM8WCEXWtu9KlOZ1K9fbz5
kfQvozIess14zx0aybW8RjvZl8HJLZmiUvzGViKaco+yrFhvd5a39O2jbVibH51tR+o+fAJ5ayre
cfJW2bQJWeDFFQoU/Jgy2oqsnupKg9XmEYODobJCR2/SQNriMOQVgMBhA6Y9mLCNwqB9AMHRO4E/
2CDYCfXebbEIVG/s5NXgf73fleQOWq/kkrt4MUCyuqw5dqTAB0jmF6eaElVDrKSdmaCGtrAZhQZ1
BP1BdRyI7jJPYtionkvqq++SC4jIyyokORhJ77cf+uxvSt9CDusXgDV2YrNggNUwcjsCpwYbC/QX
F6RunphQZnsHOW6xjfBWjou2mDwmnZOf2WQkWI9iIawdAJWapdtYBoDTTkI6XZcsgVbGja46mMhr
JGs6t2gyfdn7gxTcFxd+AzNOWCPCCsDrEZyiaR+BMv5CkO/aNTpb1ayYHqQSVhIcJNhOa59vCePr
eRlaMZtQaxZmoNLgWUVU6n2KeKhtPNZjhuj1uUWCB4todfyUiPxZXRKFR7It7CbEnhEKHIuZmnRY
c7rkWMPAvrAbQ5iNxAKeyBmhk4c5O4fx/9L2bRsQmzAQma2hLUCSQGeJY+PxueyFK012fUNSQk/g
DEXU7ZkGkaRc/O+HFVKRwCUAqPv6bFeN/IXHcOylA68L6cV3K5g9tqd0MIuetg9doL3JrxR6JBca
FId3/HKI90rTzYZ6Dv5q+J1VqI5pHgEBikgqVhzWGr3fHNydlU0QKu1tl4aLNLgYppAkVpuWmPcK
dfaXp78uAaCvPeMJW302ect+U2IGudkD/ix0mtEE4oUa6YWtD3XGwx3Z6lM7Io9y8dcutigm/2NH
JWsF+AslHiyyWzFbKg617icvSti2j5ZKI9sEQM5Fz7BIag86E1TGXurn2RdlsNmsqFK5tAUAJSL7
/UXraHq748fRDaRsamIb1oZOiQVRjC+hbcFuFwWHnkgVjrkntO7qz++FoK0xpdWRj+Ib9OMFZsK8
jrX8Z19mCD4W6EQO5BLdyQhl80Z+5zYrRqpkTyGyyS5CbYwb3h+IJLep6oVgdmKSSU1eIC2Nve1H
xr1A+VvicSXlkzeFfBWbAuuC4rfJybSmYqlGRAknsifvJWmXq8NNAEvlQYsp5YutfM9v+iPi+RMC
iXkaoDteGeEbOATpJN6AIH7pkLEcxh7I9OO+g6gOubAKYtjSi34fVlKlnDA9PS085UhhICiBF4n+
HTTXKRPmzM2js9EfvyltOu2lvEa6eYdh8exsMDDPgd9frT/FO802i7XFsEBOeI+U9GZyaQw1L4Ta
VhZNZZTrwPHSuu1mvex3AxAh3t3ESD/m1jh+q1Nt+JY0rZOw+kO1t9CJ+GnUQvlTWWXuNLmQS7Ou
dID3e4GT7hS9vw8ptsx50OzyMeWh1wqCdmBBpZ4lWcvQWonJtMZP/CjtfEs0AGeFsnvo8oR1uirf
DJsIHc/8I80cqyM8TPHsxnudhy3DHKV3p9mhvQqYebgXm6zZIrFEa1J5W2dbyTlNOGUI6pVykYu2
YnLfm6TPtjCaVOZUHzNiHSuD7+pQ0QhVV4YUjbpdspX0Fsqsm2OBt01o/C56buzEHirN7vM9lx0u
PA+qymInLMNIlmrs+FT0WwnlHQQ4eXpPIIxrJL/PZVpKfkfB56BZLfE7MXhiVwpeWcQMHyWhD0TL
Dm7+cJTfyEg84+P65Br08skMNbMv9WCyDZS9ZsorbUtP48Od/L0GcJ6NwOvsaMDe3Fihb+/2mpQL
AFuHY0zfgXBXoQ1b3f1uVNspcIwVbvTU+x/usFqJkt0EhMZci3JqfDA4jbc19M5oUw+AcDO/fD5x
itkiZrKmjQ7IA0973Jf38AcT2hmuqy0a2JssOQBZEpWMUHZHiYIGMH8LjYAF8TEmjc9+f+94vy9/
o4YCz+qDexgiU9Wv/mDVfco+Pj095xGvBwqB/C6MTQ/F11OtO9+HZ7HXzBBBInMy2XiHd5iiQZqj
hJFNeV6kR6xcONohce07tnYBe2SSTjS927sLvnPfm3wXdBYkF2zcIJqO7JvcV3mQ3JiDwGQUCOA9
chdzLaBf4SfFtIZHgyy3VvOM5wQsdk+E7rpzw8SXQdOtfFNE5HJRLoA1a3qewzJ1SEy163MxjaVI
lYx0IbDkPCvC9r+APMQBE3qb0GIntRahjK9aXQN07zxg8E2/rleWs8Fzn6UlpX2XXecCbt1+AQXG
0NQyk0aZguGpm0H53aESWDyn7MWa0pDQdWm3aWSrnzRGg7xNWmdB9GwmuZ73PJnp0Qizen+Wm6Sr
KIuIFT4jYL4i7B+ts8e9JOD35tDeIutbhLCkeLyDw4Cnpofo5YMRL07juuEXgl3xEMKS2fPMJn2r
oMRBIM8WUIiIC27Zt183/0haJo30wjgOY6MxtbYboYFqbbU02pO7quMg08bj4iNT2B2bKmqAPXhx
PSJQmwm4DPmEi5Usm3+VAoY4tLlJTAqKHfrraRIZuGJxav/GtAu0M2vz5WiOClwqWFF3kq8JNyGC
ODpQbZf+gAPLWBO/mzMr6/gYqigc+WCdLLqlDYJaoZ7OVPG8+nXCDs3lAOxFtQ3VW6pZn8OPdU+e
UKCdiQpZGce/EnsJUrSarvzta/zbsVfhMeo8UeLcTvQFrH/3MxFY1Ux8AtjlSSTQ+Ybg+qD5+y0O
JU+l0J/dZWRARTDLLy5fZdNpFu7Rij0ImXn37nwNsXYid17ksQ1Jg6PCrTp9ZyfvFUOXbDefDpeJ
F6C9LklXEnFzN/S9G1nkraD4xvD1RbnsuipNLsINXFbTodnUE1RLFmqwsZNrC//URHbILRVhZuW9
WIol63NrunJPZh2p67ZkCYdU/b/NKfJT+71UevimKUzB4+4IpUPQhsNvT0SLuXgZ0OLMuJR9TrhW
m9tf/N6+bkKazmuF5Ha6j7BHC7yvzEl8gsbKjzY7BLxn7N6locp6HdIr8Y66NGQ1JYjjwmpLpxWL
k1NO2scPEjF/gpHjSQjVBljois4OjL2SM4MiTOhLddNrxr3RsPEyyN+8XI1+zovP3G8VlAop2ZFb
G7DwEkgEw2nCtQUUAG/C3swni0pwDZraHs0XPQ0yi24mgojS10AD11iuNMnqI7X1ePEVIBLDX0Gh
aAHr3ikCbjhVObHywnML406fLpFW0noSZ5H+fIsZNHy/CkDwkejGhF6LfFqq6siQ9tPCw7mzmEi7
O2al3yEKdEiaSppYlxFcGznJ/Uw+7pzMIUTJKOSBid5iQZyU8XFC8Wa9SWe6+MKLTg0o0r6SHoxK
LwvosuJwoBdTAD67ovMzIAvf38Lyhr2RMw/ffZl7Lz66MDngF/clvK4yu1w5Fnwd0SbS2vh38E8s
/90Ulql4TWU97rhCBW9swbLloLQ9o8/0qdiTWCPiI/6E4rY6H9hpqHIl+nAa991dMtht0urtWuFe
dyx53+VS1cEmRacx+u0vqjuBmFpAR+U2tcbvVa6IStPP+LBjUBTqpl88PldEHWaX8VTD44gV23tZ
potCJFpuYhZ3Z3Gn+YM3HL5nEjGzMZSReAKkA6VKCsFsaYCenB0DMq5limSVkO1TyyrYj8vWEB1P
YteGJR3WUGqago1i47EwiuoxMSRWLcUFrHly2M9mUWE8ssMSSpFhiCsdGwvME6CdtWPyWcHuZGw6
as3cmtvYuG9wjy0bCwFh7c99SDfJPEyM9vGkg/NjrL84EnsBnoefVAO7XXwx2HVms7hzTumiS/CU
zT9cD6g9loZ01lj6qUULQkxs1achy6lzZbmUQOKakdl0nlxUxgDb6NNCNRqSOfPkoTEVfFRcR27S
TO2ZqE62B0eOMUiOkb1pH1G/v1WgO7zfNU489zrC22xEwc2WVQ982EIRieS17GdCvKoMJYqjBlfI
ob8rZX+3yoo/PZnei+mE1zcuMDcLur8g5jEQ6pWaCnHzlZpqwkF9Z10pKA8YE835gBX1L5OIQJdH
urUkoX2Ivs2yyitUOA8zE9t/F9WlSI79wCTtIV8xHheXFTsCHg6mvucTPxZ6nz0x67bjra0XJNpT
yfrtQ0Ly4GLgBgHHkyBo+ZYnxiGB+zz7UxIagY6RqApq0dtvKwSYlRH1oLglFRFgdchkjERaPksv
Y+SZ5efbQ0gl1oJozpdG3rldq1FSPWTTtu/FltEkY+jOfKSf6Oq5vBEmPDE03YwuhZgs3tg4Qvwr
EXuUjp3WYmncCjy9HPbb1G66v3cw+KwcYpkmAV6rMBMwKi/hPHkXm3WYUj9SV55t8OOrvDM0xGNt
FtysxVw985ZnkKGjtCJOiUSJz8Xv49urgF99r8+CS1tuLdCuag6+eYcE27DdF0M/54H+w+Eap32l
lJf81nMx7nIiPKxnGENuamKxC920rywHwxok2N8d2u+yotPw78ZFVtV6c4+nD7W4Ghbmt6YpnXrN
uH1yRyC4NKw+4PKbPiv7VlSiSdkOUgox8gIb8UScOi1ubvrELNIfsQglQ0/7jue9JwrGnSWepv8r
ehtRLHI6h+LoOPbOG4rt6ON6nuzCswjOvzfcVhbxUOXdgl4OV3+zAVbuV+ZtbOhRoqSfPeL392F5
Gu0h8MXNQoyr1SHcaeLzHtv/YTwWLHdMDbSdBZXb+c7r2Ob+pr1KnuklPdwcih7XbefZUyg0CH8X
JwLDfvyEHyQlG2/DCBEhfS+NFIZ4jcVVdNP8gWKThb5DXQB4/mtwaBMy0dFubfRJocfq5Kl5LTsP
gO0mIx3JsKMz02PWo0oatSBa2FeUeivclE9x5ml55qMU1h3d0Q4worQqL6a0uNuiR28q2bkgMg8Z
zLqY9hoqI1LD+lrBEm/9aoeYHUCjwvGzwQqvXX7FoyRAd0wammn+uNLk4TmBfMwhW7uuXapowUQh
fUau7QK79Qk/+ijN0zHlVl6cpvgpNv4qTo4cnsTa2yFNaC+eXwc1eF8YWCjKq5hxHpDe9Zuo8ncR
57xtN+IFkF4iEmEViSVhJLzVf3oOvsSae8VjNEybBpbaQLPwtBvAuflcka7Nco0lSbgpxuA8/yu9
KhL9F6OqgPk0rv43v3+VofP2NfnECbYhsv0irSgbDE8nO5kqU7I0r/t17TuCgvnm1g2sFxeuc2SF
bTh69f9GFu+sRK8knwIYfFyNpM1Vua1bALbwJt8w97D9CkTdbssGmmefdIl0RNbgrvpYoCWKbWYd
an+MP4axms/zp136SLzx0lAtSZn2hPUHs15ODbe4yZyQ03LuaQYOoYxRFXMmOcEj5vBoAw3iKvRv
iaQ9kU8KBj6Dczcm56uZf5fGSRnm2RTjZpMOA/LdN5kQP7Pvy90Mw6cCN52qAh8AdYJUkg0OvFoj
Fjmtx4/WiMcNQqfnStsytQWhUrxODcO1ywNTGtjhFHM8kra9ABSp0YsL/rirCQPUrmbtKLitJ+Y7
WgSXcqFdOuWeQQypeleHlDprE6n/6zkowIoaGxXOy7KEVtZ4BkeYf95t7LU1wyb5caPo2afQW15U
ZS1i5C4t6D3rK+GgSvLe7Gadrq5aj9wu3TZwbfaMs4/RCnwa2izqqhA3a7TWmVkVD1UNqB+NCrWy
dINgOhivNevsFnljPQQyVbjrVu/TVeggq5U62oCPM+MLZKmx5HZfwM+TAGfySF72mPEHMNtcRryJ
GSelIOg6j97Ev2RqmFXkYZa+Aw9se9CeEOp4XYZSK+7fYWli9gmqISdUrdvjbM9RRKK4ZoQ6s0wG
lILUj1g9Nm6NiMOSwh+R9/2pq947iw3xywjr5oVAyFohGxEpD/Bq55Pc5RioaUIPnBpCiOyW/6wZ
OF8uHJ5Osd1oWNlUat939m2nMBKBqIMrO9l0RQ2QyVoaFBmaLLjSlOTqcyoy8n1++TsDAmKa7S7h
ZTD5zQl9C0vBVhfYNkUQWXvanx52mU5u5ilu0tOI8ZCag869HCSwjrHbfELHVU3cUNNsM3x3eUjw
dVfPM3mGWYXFy+nxEdXQZmgT7C9Yncufq6wUwU7TQIln35oKMdAszZ8Z2DpW1AV8vjH5TOntbfc1
OVX2r1Jlo6fsuDeXWJJcyJD6xOG3I8fdkaIHnORoAqZXBkyMjzUpjNZg5mlXYNVpC75oY7ax1RyU
1b1A/BEH2VS3soC4lUR1zIpne3zunarXCtC9CkBcQpQnEX7aZ+MahEAeNVenmqkayUPxYl1JzehR
sSObHhYC2mSTpv4+Bf1np1SBsB1B6Z9pC4Bel930sWEiTebZ4ogZmwlt+riJC9TJOM1IPynm2ckC
2jDTkQ2aoimmJWqzu6MLChUmmHgNWntN2ARP1qhyuqecbRmW03AntfNRP9CxoeQvadqrqxiJHFoM
zuVSg63f7uG4sVf0+CYiS9/Nc32+Qo01GxbSgLAy2JWzoJqgoiIHGnRUo+o11uHq2vLNBEAv4QMD
l9UIl/QujIs9Oui20hJZqrD+tYK4iqYMZuyFTzimYvaEyiU2No0Mgxe4KPJcz1YOAvN2deCWGzLe
ha6MBjoBw7lElcsbZMHh02QJqLQ9HdozjDzUdG0Nw/4DghxpuOSTt+2VVBWdHX9K/BiAjnKLsyBd
1hYgm74hM+UDCi6yvfBqIu/+l7BX+xxOrJuYg47xSPES3BcZIHx5SHagUD2swhBPMFRs2E/83O76
o9xI1C9fa9LaA7fqQjZRS/eHXAP0UnEqWREATihycBJ7Rfp1SVh7zWmOXIpp+mJG2tIC0ZiXjkSu
9uYlwyp5vXxzA5nxWsL76WT1r9J8bFXNbHKr0Sww8jxSiPKW3b40kZrTuP1aUefrlVkgKeWjSBhO
r1V0BNzKSkNtPYPPL4ijvtDWJxfYRSqGM+AALUT1dxazm4Wf40bSe5R50H9749SosNwj25mifvPO
+wMmbVpRRCYGPz613CWNxqqX07HUSQ24L+GzqtXBY+VwzK7gX4spQTmBZMc6dEteF1UhO8vJvqMb
QaRPSqMwtJ4oM553Gk0chYj/xf7V9Dz2bzl7DdSlAmpTQUP/D+03w2sKAuazzck31E2zURnSNSw8
1VazMbfUxkGl89+ndHx3Ha1TSsAdRmUnhfT4VQJak5u0loMR0DjnDYlHtVUMZT+Zit/eNpFuATt1
kpIkDJlLWCz0E5iNTmNBfIof+hj2zlH1v75w81az3K6OvuKtpam1JlzydtSf+zUyAcRLsRXm6HGH
qW+HO/2VZ7yTeJrAPtYSfF4U8Cts8nLzbCk/lz+hf9uIe8d7aokB986OvYH2XsskK8qWnUzFnN+J
xz2doxWwn9A+aGh00LcByc7LZmMtQXTzGz8cy1gS+8dXyeniZoFDERYFBPjMfYSqsUnG3oiB5ps7
UBlhiNyIPMILO7JeSWXMgiGJdCKEo4XoN14+WJkNS9C6qT+I4Xznl08S5k3VMsygs74ydtY3IhET
0U+ri4PsfPMkFRMZvtDNoDB3W1vhXE/JWwF2b7k/8hiEieLcFccwsqPN+viPrJjs404iXKhvua1m
y88MnNPaYqJxxc+ih3z3dQEZ09eLRvu0B3yk2w7/a0i/lnYmxWt3aOlmwejIydQ2MDkGiOO+iURO
Qrwo4/Gcg7Zd3/ljbc7ucUonEtPRfzjOBHilA8YdGxMxq9zfC5WF/42SOs+aMhGxKIUklAjhzi7z
KL6jwLjWMcaWI+Gsoby+UxYtAObUN3vAbGU5XA0oJsDrU3YZUQzSlhOohrOqFXqMMYKTj3FpG/BW
vmgCqLW5ITRtFyQBj8iXDnQ/lzHekboecPLc1gx5MFSVJ6j1cn0WbRr+G11fYAnYnfVsV1Onlf4N
/kuEC+0+VBHg+T5IUeUHtoiJF5kb//hlZwpo/Mnp0ab3uIQjISbPk7Z2IjDCSemhhbSkWkmYIqZ1
hZVkoJ9w4i2RgHQfYPUj7itkoS4FOm66KiB560qbz66c47Iy7qw+BwYd7MW5wG1Wckw9PD90+RnP
1vkpjZlZRe8TI4ysqGKJ7d7dVRwXHH6nFobULuFlxbpmryrtkXJF3ZoCA6DJtWOOsR5ugjrjCjVn
GT9ozKYflBOK0w1sTE3EmzXOgR9DnTRfA+Z1LH7qqA+RADl7g4kYOPE3RRiJOSW+zRu+4N9VsRZi
vt/e73D4OjbTkvmWYulZHc1bd/DJZEiOZzN421643F9tIIcpZFOFen1Yd0SSfvYj40VWLiA0lgSR
ucANb7AN8uuZ8O17EGho8AMP+bq2JP2XqfoKImdGDKiQ1ez/G0s2eW0wO3i70hkJlWbRtJpDJLX4
vAmIMebgil06Dukpqy8qEXErieb/wYzuB5Kjs5iCSmUx6vBRUuX7gngRmYotx1GCxMpHMQnx2egK
CmgCfxouhWMTsZz+WBpVS9sr2H+StzwuLQECwcFmeGap/Gz1htf68Kl2bGVVQJFERNFYxPmtW+s9
3biHUrjIgnEvLhCC7eBjpsZGwBwd/qUKTadyb2yBYl1HOzdbhepY1Nkfi843bhA27DGvt+Tm9Xyp
8vibBwddzyottXpbHukQScaA5Uaw1PlIZK14u7MphY1Gk4fpW6LwnhwNHaawg1CGV640X8acSOkB
0bavGkNQPqzdLFOoDrHe8MTLPFTKEpiBuL7KLGjpN1Y8EEKl7T72vi7tu2iuQ9CnuvdiKuJIO6qJ
PORLRJdM0rxHyqtVX2bqcR5XQDX1ljStw7Uu2AUBhasgnaLkZDwzgSlGjVC0ExdGL+QN2iNGF58S
DGyWMB0Gy6WW48YtKephppYPWJIG4cNT8Wi0tVHVAmXp77w9GhCme+9fblMQZG0O6vlmTZtVlmGB
DSJtxlakPnwthghmA0GXtY2Qy6K997xH+uhvokaLhOeQ90hrd50T0LdgJIGz+iWbhHuhxts8X+Ru
wG87uqMl9xgYi9asVP58knJvibQ944ViYDmmEeYFeM/c+9xePla/qTcbEaGqY39FqGUbH3Lom4+H
Zh7EHUR26QOxozICGf/F9+ycRoHKS9bNoOeM69SrROfC7ocJes+P3dRXxlzxq+o+46OKXMv1yVU3
qbjGBfDzdFDz8CKLDVRf4S8ardjd/Anf+Vb8qEhgJajfPg+GI4vfJMhtD6lbriPjzjybtoe2g3u6
54zZGUnTL6r/TMLSOX7DS+qC6yuIJcPYMpdSKA76Qbp96Fw4MYqO0uQhyPkuHrzv6LEtOMzrpzn4
QkIvq1SF0SrGCGTPdKsLMzh2yklPZe37MV5f/LaymqG4q75VdOnMO2pE9M6la1Rhz/Aftx8YvbAU
MLG5XtnH9MBH5Ukf1mXegp3wKjzNGFiO8ty/iPrJXYCJOFU4cJsypNDE1qPJY2Bu/CGoEd9DXvSs
4dMFt9MVvR6lmRsVzf7Tpv6aO9bRA9Ambfc7Hy58C41gRf2+3Kxl6+1TtvTeit/1LcaFyjxaBCO9
z//VVEtY++jPRFYKCTJZfs0O5gut+8OsDCIw9QUiJvKezX1cAqrjboYlDFRjGL4KT/xOegvNktQv
lAEaPEvUp3nP0JhsfjPavEcqxoDkDB3EcCcObhg8q8SkOtUgV8v3WWsJa+Huq9q09KNzPYiB8sZw
zmwQhQkt4g4atV1TFv9i1VFpj2+ELH6xU4FXxmO30G8nOAU1yg5LyqpiTZuWANJOpjJVDrxynQZ6
5JUFqz0Iw4C1wOFGDvU2UmA/Vc9+nLNIXnUEyrEV5qFPRQm0majc8cTcojmQZYuEihgygOij1KiA
rNpPk9SxZsKu9Ovg89OGqvargNrVKpxML0UbMBaL+bfh4U2kvdrPWkWxN06hOvbDboX9rosqyHS4
nv07RYkQ6PU0XCCggC/ruydNK1gcPteiHaOntPZkQkZU0a1pY7WQuu7b7mjY39WXDP8pdFwe+V1N
AdWPZKD8E+BAzvGFTJgqIe6DHdfVc3yX1nJsNmuRELugRl4hNEGfeUkwfLSNhLYyULh2+iSwm2T/
2sks44hLsGhAkcHWDYWerJn+Gu+UTVB7IQ7eonnICJSm0THl07RnUeW3rI9UIAQt+JW0dsGa6qp8
AoH4aLhzruj8OomhfrUn55RITJEPVDq3f2JMifBaxFeTDu0toWWSiYng0nNxYO9+a31sygL6vdCk
OpqTlsZ3g2s33iZR8y/+nb1P6xVyR2CUN9dYpTk10rC0A+DgMIV5BxmtnDT4VppSQNyFm0l1kLgc
+Lxs1x4xBV0+FKA1CYyStpFB/XCFq+h9xut/fIQVEjepgT7JmQ0gTBuTswBUFNBY4vmv/VgWwtwN
tRqlUueGWZ57ZUw49aq3nvb4n+ujPID5es6R+pjmeUZQrl99IMqT002tu9NAhPC4RQINMXrP7mto
CL6o6T3crI4E9xFG0jxeysULDfFPPe5T95M7BWyI21WDXbRjnInmPBLbhd/u3ySySV+C6aLzgUvb
NTPK4Gm/YN0ABo4gF0knCEgYzoyVamEBoqus4BySKZymduoZb2HKJy1zpvHVavLyGq46w88aX7Hj
p/dxlp+Am+ESaI5WpAR6sZu4JoRleQ2ITnehH9OVxMij8v6IBOHYo5OR15PYK+35WyjUXNZmX8TC
zpwsImu7WoAoNdTzT5k5qLEjkM1Fz+E5k80lLSlYt8burv/UckmcvFdfulzGAUb03id1hAvNSgZ8
Fbkg9C+fw7Q2mFTCEFGGSzC2QSv1XwEJe03JMUvA4cr7YmjgVRNidMlaAcmfoDIKbzQnq08nqWVl
NsXx+baUZGFPEjb0oiTQJADU/ZMyTaaF1/VCCUjzfp5EoCbAwFc80iPe2lQPFQvkzpoPVnp78fT6
HW2EK05UFfWo2Ncgq0fOSU8bMDLzIqPO5IEOnRBXn+3xIMCLcgNwnUzhEng1eNJ/ybsKV6HTU5If
7pAX5TDy5uyTE5+uviAeA/LH1wIPiKrvYfroveYYpegi7KPjgh56pHIsUfv6783cLvr+KB+CwLx8
sVYXyIzeMLNfexyhktH7rlZeYzfFBHnrQGtCSYZYY/RhtUaiDzjtNAcftgulXBeManDTEA0EDkJz
CCiHvasJCWZmn9Kh6uw4IDNumw23TTY4uaIkjzOKPn3dh5TxAtFDrmTgZjTzFQExlSlQUCQwgJio
yKwNl8OgzRj4E6zGsBg9LVH5g32YIfNAWLhVGmSv24q2oP4kHAM0qHPG8uO45PWuxw3CiBEPnRbN
IqtCLq/OEJK9FOpAwj+PmAjzf3OutJ3fPKDp6H5IEQus7FlU76Eqb5Gqlugck3fgMtsC438FuDfU
k+77CRHLZO/yjynwirENSQ9A2xkZdkspOOkg3Y5S5iAR1V1UolAgmGu7/mPNkhEicNaaW9gwOXvn
fVXrUj4SJeThm2Uauwqqu9YrOmC1JAT9gcz44txNusEAXrhte5+h3qXtIaz7iyn+MnFLprI7uKy/
39aaDVDbrgyhR1MaW/5dpAZHu/Z380ywADVlRue9ppDGMo8kid3uJhsk3sekjM0BhjV7tT4DnCjc
7O0Cod9LVz//SCbRYITZXvRVrLzTjjwtKSfwqDuM5qQk+koCwVlANiDZLCtzQ7uP9Yo3AyOVtt5Y
SsNA7Wd3V+aiYnBaI79l+sbObKEoi3Ex5YCD0TZhK1+3fYMdxYUseqeWDc+avQ3lU5PwqiccUfzu
4hMdd5SynAL0ekYKbygJlllgDdOY/6KrOHgWEBB6xVcyHZlJ6qeahj2iByzdeb8hQ6oIUydhPMt1
uxLWzcBq23rIeO7Md/63K5Mu7r0EmucBEAGOmv0F+djLhbYS2TsHrO4AaiPT1I1f2PytcD7l7sbP
curnsJr7MFnE92AAiWQQh365o8ygVWa3qrl0qzGKKvEGagzCD/9U4jdsra49o6YwboWjZpxPHMi2
rAF7RnAkj2gdTAaZFIc4lIR3diezK6CEY/75AJI4wfLu3fYeUE0OQYBnSKPpvn7/C6nlQgybR63B
s0sCFSsHoXgLL9NgS7gn540CYVKgCamOfCL27rfOyS3V0HwBJajepizYnKKNibWi8Dr87kPP1QHQ
Rovl5rh9eC/KaS5C4JHWZkMnroJ5v+Wq8gnreLnt3d0EI9zvNk4PgmZGhqZJFujJwlHiDG/HnzjQ
tl6DU4XXsO5haaj1IP2oc5/QfvJRs0ZrX1t5HeoTwlm9mbou7Q/hMpuR0S8ItKM67ABOMGXiOUsa
/zwy4o908oLY+4Mszo6OxRFbnvWZ7CG7ui6W8YoF76rgJnUqcptYNEPUkRvmI88+dyMSfc1DGcnr
fLuM8Ul5l3DVXIgE4/HyDZxEjFJ8ai2CpE5PltwjvbgQNGWynCRtJas5uB8CizKbksCPpdbN7i1o
VLP4wMMU4sA1fEDgdiOAJN7Jdfa88awFZAFoqqsCl5L5k4rUZxL5o9u/dIC+M2cqnxnjZWCauUQ7
iWtz23ltoDajc1PGwksgkIH7bqpi8CR33AXDJ/0SCEUCn0GPTTPReYr9hsc5lx1wN6E41+QZVtRg
ErFJVF7lEGfBEDk3dDEuVovd/GaYiwtWObVO2WFTJ7c0eyDf6veKoKJbidJkonbQ6KlpWrEAkocg
XOqx87zOsGjEfbiJ77haSMdhoIwRn8d4Hu/ErveRGA0QTEDMg5yIoF/bhWta043rBpNk8aWX3r2D
rmW+PUiHXOX0wqBAu3BmAGiShloU29/DBGH6/tR1OrrzaGxZsIoy2n4f0rAGANLHcsVHm9Q2dLbc
LyY+YoDlNxUeJdhh3KZFmmjyk8/VzPgk6NS2xLM9UxakIQjSEt3xo1BNHGo84r9SN4byNQcA1NUf
7qK2Lxtnj5wqNKQ8NWw0jrhULE9eJLsz1I7CPhfkHFjIycccI631EL4q/BZAJlJEW7izkDbveyPN
J8rdSBrLepUjqvXEuhEeHIh/LsECIxMIqjFULR9hKMCf2gH9PtK4IxUSo6npxnpYn8Ihg54kOgcm
dAAaaYfAAYepyQwoU/Zzy4k46qNy3we4C3u+W11YA7UXNd/sor4Ki1pyD2mN3qTlbsgTBrnIKlFH
qDeSEaApKJXKLFb8F8sb/u5ffp0BYoLLrYfYd9JiP3YEB5wj38W/2UBzS4xY5aRwDkEPLNRzKzuK
w2p+kgYkw/9K7X3HHqU/PxJbELhO4jU5IpVJOta4NjsQ8f+POynRdscE0XHBYxC4v9jFvGjrHgZr
Zn4/WYw1GdxGzmH04J6pHk8h5UQwSFghxjfy7VaatXm1O4uEF5wUadXu35dvIcGdgJ5oxR1GomRs
r+M531pF5U4jP1nApkOrurSFCDqIJyUVSC85wqSSl5ULVXlcrTwdEGaDxu275+1hlkJj5XcSCEX2
Awj+Ev8JxMBAmY0i5FqC3r5Vk0t08WFXcWM1vuKYoD0oxbS7SuKxa8TalKtV/BbWb9nZyFXV2Jbj
w2pQmr96TsuXJtM5Cb+T8mEC4q+p5Mz73PDgWrx7VUYngqLR/VMh2NaPPPbbrqYUTRT/xn9CwM42
WRy9r4zVx6usM4/QQ9+/4qdXvPz4phSCy2C1eWWmW7wZAppSumcL2UTg8SxytFa7RYQuNDtLyF+g
WUc4iwh07gQi1YT0YyOev+PtxRr1pefiST+UywGNxGPhdMhx4A4yRL7j+gNErkib7Cjl/jF5UPxl
Ns5CNn6JlVCt1UDoqbSS/l1+v3iJAts3N1vjmG/l6L5/g2ddbhGQ6euy6YwuOBXkZlIlt3REboju
r7TFyI3RGGFCIvItelhwp/Ernwn+ZfPIZdZy+P1wpqNsguv5ECjMN4bJ39xYSUkjSkEjOhT/Tl2B
vJTDy2xXN8tWAhyI0ySpv3dE2khMEbg5IpKYUFd2vEJRFD29YAC0W/GnQuvMMZ6p6ZEtSFA784Di
J0jKC+rMHQt21c4tpaWXngRtcMBq6N5DEVgdLJxVFfAgeSK9OJhrbuf/ZIhtjk2mPXR/aW8rHjDk
c9GCPy6MMWiDDTHyc6J2bkX+x//P6nCqk/OSzCwIVhyDhJMwx4AxI6I5zE13gd2wFVrHl0SylbaX
d4fPPuuTWmgKt+jwUns3fvlaecnNob/AqLp/Nn6zzdKH1JwCDAbxcCU1pMvSBVKyNla4NYKdRPDC
weUMETazvYEz0QOYwR1Qeog1NsebD7QiR9b1TxtLpg6/zsG+4BdhtrGyJJXtLDfuOs0l+yMRe3bM
+AS7sF14ZrJfZ3sEHRSZgEXvSq8wl2EKmnNnUUFsZyVjtc+Gv2h3D5leEj9MfVnxZdiFlYopSzdP
b2G8AxPB6Xvj1oSE6iNe06XfIBrH+3uKyPia3xgQXm3NjZkoRzYu6NPYCqbjAvddbFJS0aC2sGe2
mnlZRSjMYPapZhxChyfIBJi6ePBPwP1hvk3wjZY4S8LI3xqD+ESLJlZoQ16qSzWcdSm/fjpEnNCa
ZfmzYZ1MHm3O8O/Zf4SwPhliGqpHRDA+7fMS+OXuZ5vkdml0tYedc6nqiS5ullkS0g8yHndYYqcC
Z4rm2thhvskTPKYssdAmIwfM7HsROEV21K4jpLVLz5IrMYMmv9Sv/uF0vBqiWbISyZyxFZvjLOps
bsuCVq5xgh0puj6tgDBdAQyj49N6U5qgCFu1dZdUt9lTwsBPtJqvcj70zl2UGisvRwjCjgONv9Mi
41C63l54NRzegsxyEyMkNklRBvhCZGtOYJo8vcdg8FkUE3mtWZx9E/weR7BmxW/UT1OlqF6nemqH
ExPP3YYbbO8R6O4B3U82RDynchqq+5lnUIm71PEdJeD7NA1ibkuNY3Mm6nmEoIj4jkJY76f9xR2n
LhNX5vwNb+CaKSNqzdhrr6KzFMzdmC7LaDbd7VxJFRfDqKz6bimfM5FdfzcXbCbwYfEceQh8fmWa
ECueObDA3q3K62wumMj6HMuYfyJ0NbpjZb5YFVDrL1a6TdyLDhFWn6NKzbdwcBKiiOQdCxJDad3d
yP+7SXBhBTyGeHDYnh6MUkmfeD99J2sAPicitY9jNgi1jwl4wQtjzCC9K0KRjkzWW8fNUlJ9lJRE
MqBVuQ4J8R5jMguiRU/z0QGESCR+o+hyepnX/7qayEq5KzDV6ix9MvrDmCrkD7EhLcX6V8dL9mgC
WdDJ613o0DAUEj40o/Oq1Z/T2vJ1c9xyGUC0zr06RGHdlt31t/XYMxvB8Y9jLXIJGBi2I1bGX7pN
XKrSjvq3oec0Mis2wK4OpPwPbXSPnuTBYBSNzBO25K2fdXwf41LgHa9ZH9x96UcJrdpBKVHjudPB
3YaJgia52y0lmYBFWID4T7O3J6BkURFM2gJ+CpfePJbNrw5NVgxBSFha+LTrJIIqBVM9iWt+rkZu
M/4fWDUL8mIxhFIHhfq0K4Vu+eyn+pr5aZbMm7Lg1M+IlMXz95N3Z17RiZRkMTIzXVShFzXrZJyn
kbbFOYH1dbamuFiMQZcan8CW1Rb+iDIUyFFZRfbSCsyQ7I44PwUcSrBqW02EIz0wo60ij8KLMAXA
2zwLngAmOSSVo3OqQsa0Mvd0ITJdarmY/O93+aKXf/xs56pFft/14E8NKx/aueVqCdilufn+valA
LrEMPCZn6Qlv05ylT7gh3TgXziuDkn5iIvJ91CK8akjSmJIa95QlvU3qlhhNRA2U4N8Ne+NNobP7
Di+RFU1VCDAnj4h13+VxglRVudRge769PYKAYJKLfvf5ETqOXg487Pb28L1MXpZlRcf/QrcNh5Yj
utnTppoRQtK7E45slEC+cOA1jYYTwF1sySO1yQ5bSOxm9UUSs2WHAOvQXEoNqKPOXdrxzZsXMPoo
EP72OoWy3fxhM5Ds/jwzYK+tXhL2Y5uKvIenPgnAsgAvtqyqgcMhcPACkOMj9NLQJPE/zimIapdt
D3ASCLkiRTqAMu2spgCVzOJIo+Upqb6L3RtFukq2B6oD0sSHrxKJK97tJX4dIeFeS4hKXOhPM8RU
0/qL6rCq2gaUXKz4geGlOhsyAtTPsVFelp1LJ+ERa2lyas1jeaCYluoaeJ058OkK8V9KHp0l/i2O
McHpTbn+Fn+7CGL1ySBi3fdA3Z51wHEFSOXjZsPuSdzh7JCrsKkN/pm7XxU1aRMDGElxMR/aJ34E
MHfRr70Ls9lK8zcjeePsuILzxo/3+rUdxhdZX28NNERiqH62g/B3iNfsivL5XMO2z5nB+uoNHjl8
rHt4w33R3CzMDd+bNFK0m5tZe4/FLjnNiHkK+pnkvpuTiYe53NbASgZoXjwtLKCXSzttSFwciZKf
jdcQeaKUI9qUKmmwr1KvWO7Y84n0ww6k/2s7lpOaS/nWPUMU8BKzcKl34KEz6iM5TTqq/3pMVgO5
ytcfKRa297QXWnuOSzMZSULVFWVLdDsBMHYkszaZLHVZ8qNRFmg30ntSPjyoz9AFThCe+em9lkZz
ttZV0dJ8q69gpuAnoB4TKQmzTtSiRCXmgEerY8PDTw4DZC0oX2AZOQKjhlB3YtVYE9JFmOwDAoua
eaUa4Q2xRF6kTw02LzzDU7Lr4CmfozVD8C6y2X/JfN9hZXlIVdEpOkhJb78SeQooHUfj2oV/eerN
z9RZyLH0ySsBrDSMwAqxy3x67uz9/IHXFdThy4FXPKym/9mo9J/PEit325UmlSi93KEbxJ9xrQbm
0QbODqj40SIKiCns9IQiBHbuC8JPF1ZV/YXOGa4OGBF6F9wHBc5sJqQqFBrL0rRmphl8rDSCIjSu
9ktMvzr/yUnSyw2KoZ1YYgrSFXYvXBOvBWFj0MO+UZl+a+NHvio48nKEqzH8bXHDapyBYTwpzeAc
aAt8RXsIZvc5gKS21g7ngyyP8qsrcqceZpZHyKwwKhyYYDvbUnwOf6gMxB2y1mNtL1pxvZZtzao6
OLxuMe2xMZkQOHVaVTRTK+xtZKBiUg9r3cF1Yes6GhwEM43EtLvr/kDBBu7wejt0pYj6ARXyev7/
8eDrZmiudtryagv913f2DbYPkqSdgTbFC3KUAxC5i2UXSaI+1sL14SQQJTuhMgCbaX+5LpB6o/V8
Fm6vNDWjJEiDy2UpyPhHrDjOtsGwFdaUQHxHcxbmjjFCNqAviKhoUkhujbtd6qMdTp/9LdERgyvl
TxYs0IVWWgWlYUuAyknPxF7g1VuefbVGAXIFTB8MEoNUGyImmASV1uSNQkuRG+PPsJpRFWkEo9My
3MiElA7E17ZX9Ko3cfwb1y+Cc+MZH7X81/B5Obt9BRynJul9pq1anpl6QZwEl7coxSCHEIazF3Zo
0jhftkDwu8zWUsx1mrxQsrS8FIqAnHUBojJFps2ODftkDFXFGRi7nsIb2z9ZQylpkZDVr/UxBm04
SLlVAiD/CMw1Yo+8XpnTmUyreBWF8XBzBaVIFCBsL711AXKkXn6Hslklkl2HFgalSnFKQqEP/+ck
tnsmIXCU188pLkwOku45WobH5WJcejruirvVFbGNkk4o7tU62x3+IlxjiVgJQ6CEFcR+4K3E5Kki
sEnk4VPPJxgmVv3BYp3no7X0wVa1CrGgWmW3H6ugDsZfi0NHmDeMz66lPh7IpD6GwvVfXY5jwFvO
uuoeNTNXzJEMdzc3jJfn1N72+2JayoJsZo2jMAnWkyPzdPv+T2XTQI2vxd7MK3/3mu+jbvnKtK4Z
6m5OWJkhrckq8VsViKzyFwOfJKfuio8HtaGvTDNn0eq0a03DOCVWPK9hYDc2snYhf/N2AgZxIIiD
zTQLm+XoEh8zClX5YjaosX4bZiljc9LYKqm3wSikJ3DrbyqvpFDO/kRN+g7MKC/cDDVexYnBPQ2g
I7m52QYLDOZhCZ39z4EUF4Izcy2eeGW2tCB1UIMNTNfF2fsL4N876GxSPb5HLjdNpKkOEnrRfCxj
nXpU/SqxBePT66pkjVdvV6qPnzss4KZTFK2jDScOe77mcqFeazAfqrPQEidlEGDUcVc6CmCabA3C
e4XyCVtA+sHYUB4JVS1qCaau9JvcAutQqH98CoJHqsY9O7EYedKxggNQ6lXeFpWaktaIQFnvVWrX
XHoVpHLLlWhLTVxRvHlYX/t7JG7EI6x4JMHSuvYIXJIx+ZNkRc26zTL40B9a/uHPDNF3qqIZ+8XF
Sb6NRQc0WKHvlFJsoKhgU+JRSgFO0azwW8lQXc30F1cz7qCUpLR+TXcPaTRzqPcTFVVnILsAEHRr
l/iDhPDWC/wWonXzQdmHDxZYoemYUp622weRscmg716mJg7dhjHzcTT7wgKaG3kh5ajqJNa3xDD5
9lpSZXm007Rr9AmC8tE5/1W1Kb1yP22s5XFDgCcqjN/YKnBLlTUAay3qre4OwUG6bIK+/FyLTFWT
qf/7mQJBubTHVD87B1ukOwFUV812hIAF+dm5V5KZIyFxaeRevR34tCIb7rTy64vkWA+dj17kuwtR
t+cHyaDu4jgsGSy42mx3qUJIeBTb3VUg8IpVTdAWM0Uk6o61Nh9L+93IDtrxGUcrWPrAiCpzKtT2
5HP44D1TdFcDpdgc3oQSSJBy7Krq/9EEsjwBF1sPuJkmNZfattorUwC2PaDRIBdqhC6FeifGsIPQ
hm7dkAlsY7wQ80fHmLnPPkBPLu91yj8RjMj869tG/SGKICRdjUR36LqXxiLLAFKM94j1MSlr3xKC
fZ/PQ+jiGZh6Cl6Vs1QsZVaTfHei6PL+sQOUfpmwqkO86Jaf7VpD8aJ3thQ0BOQN37q6/94Kdl6N
gbWIgo8PQFyPM86FdXaAG1hN7qMiEXNPRWRAqinCkAtnfwQGF4+y4HatvsRxsxqgxeeDfLiqgoX8
jgFGaLabCrVEERKzReuACdgMOd6n5OdQQHCAuUIKRRw3ZeXpCh9HBXCVIHQ5MhhPGNC6gczUQ5oA
sSxZKaxwZtgr0Md84lrl3CPEo/KJ8yixGY+AxcQFlqK7/HOpVHXfZO0Bmf+miThR71BaaTgm9fv9
zbAkqBjdlMjHVe5MjMIlWrlJuWD9WqnnpbA5LISMnhHgMw0eHQvimQKhCkF4MTgHjYNrTOzclOTs
O3CeYoZFpnrvzch49rOV79jYhfbEcpFF8KE/ZjsNfI0pwXw4WaqoMJ++wU+OXHltw265MxY1IXhZ
YliCMZssIOcBr2khn9h3X57VkGiA5oe1M8FNaSuuDEzKEOefUyOYAZAVBz/uUOO9EM+6xdCWyvTJ
jBrVcXO0+WJMJ0ccaIdImmqcNL/tpgT595Zd5vn7Al55Ncj5zXCMYxXCG+GgNcPQvk/eeNOz220G
S5B5b6z3v9dgLKrXF2VpU+Rjl4BD9w45grxoH524qEyqCbm8iCJzGVFDzZkK8mt5t8pQXn9bbHpU
3jUdfGAf0Qjjv2oYJKKUnxnbhTnWKnr64V5D7DHhu64cuOIwgammWGV32xTseUSkuRmTIpQAsIck
Sd8R8tjTnSr8+odrubsrPHNhyiOz6iTfDSc37yDjy6M1+itg29NHULGgLnuNdlNCSDrRiPN2RkOk
3HwEnU5bw0WBkY8fmXRRkfGHfDFP5EQaFrJKSdiW4ZlDSa8GBShs9oc6b3t1AyLiPwlOKKx9VHDD
0cU+oAWiD6pxDWq28i9KskhHsOrulx8Nq+XQYANTsAbUtQDdr7za2ZuNQP0WbXruIZyODRiCeRVy
NOURjjoHnWztPgUyLYmH73wyh5+4IA2K6Ek+gaKL9uGL76fjika2rr8P2HpcoAHNZBkA7jQYKviv
29folI9qvKRn3pjAU6oLBMWQT3m5z0ti2ZMV02lRyLRtto2eOwcA/Oz+j3m6/CpK7AqngFFkHqsq
nA0ItxKp+Rtd+E8vtphwIu/+8yeEwoeTXpOSkUWqq7uJPVjHo5jPACFctb3Kk+ylB24tSaUBuBKL
gVNqtWpjzZ6WtwpDJVFgxYP7Yl7R6gj85GEUkkF5qMiyosUbo6/dLORH8E4hmStFWpVCf4G67Ehc
uF63B4i3jyj1Eshr0HvgmR+GiomWvRuEa3/ZiZW79KM3Bo9sjhvE2TXYbU1Rfkwo5dfqd0CRYb9U
h4y7LSg3py4gtfFSCAXfINV9gfaV0Sb1xkrzvtbKdaWXh/gI/RDkVEX45G+FKzzDzzyB6he+g4D+
E5JJa8W2Qx3HryYwe6IuDYDGWtz5sV9zI+YQgrpBmJ4dwNc3ALimcQb9Pg0AHwqfYwrskaSKJU4V
vS/AFqwHhD2Zchd/kAj1mrVdrpx+9K7C9YfDqHjIUFkvgr9lONjcmsFOBVU3z9qQGAFlQeJOJwWi
HVZ66rVN0wKENJKASx/khoTyi9i9ahQizuvqwcnAsj2lJS9s11z3ExgYGYMTOsusTyBVkWjTeVlP
FGFJWil+7Wj3HRZ/8Nhu/IfZckguFErEsvIzUTClC6+Y7uyo99vI6YfuqHw/6ajJ9T3Pe+IgiH1n
W41H2nAl+Ynq7g/rGeN38yoIG80aS0XrAT1kFxoglHR9GC6KJ811TeOfa2zxEKoTikgJKmPVbN0V
pKz40ab/MSgOwh0PH3lCeTPt79MAIaEysSQdgIr1XCF6VCVL4UjOePRo2c2OOqu+uBhRshSYNZ1a
Vxo8fnsbWQ7yqfUnWGCfGrrj7X7YBM1GW0KgFVUrx1hp3mSpc0VQ0m4WfrTN6XWPmIZFftE7E/+Y
rnayq+FGT/0Y4ffuHnKEmYLV5mniH1cv2NE96QCS4R+NTgJFLAhia++x+XgH/JNRMUXUdmm7pveS
+uTSBqKLgEaydTL8Vyy8Urckl9evYHbY7hucvTUH+vw4VtmtCUrNGubBoA489NW92gNhnaic5IXY
eK+Q3STorsDLC6QV7otwtyP7oPGVEfDUgAxcUwhcWh0jXbIkahFQ5g8xj5AOs2Yntx/i75gJYsad
Bqffk5y744hxCiBkPJjHE6wF/yAU0p745zp4T9ZCIKp8I5zDKyeqRNBeOUuTIrGZFtJS4KzPODhr
cikw1PO4SPUa8+25HWpdoLNj4Uj8lMev5OGEWrCovHFkCOKsJxgqV2Yd5W0MrDc+6AHb/oV88wld
alJRUeP9nQcGl6IBEBR7I8su6xyJJc4WDMx2XiDXPEMHa+jVj4Q/4M6SdKJPe2WITwAA05YLj7FU
T0oRpZvwLOvldoYQN6R76uqEaE3W0hZmCM/IH5fuE8dQrVAx9fP4ABsu0euF0lN3jca3hmsfrPqg
m88BnGmYkzM+E3RLkq9OY0Cx9d+9UxSWeAnXejazzPYCznJJaNJEuDz0641QZjla0VJutFMcAKv6
Ro88OjXKzMoVhcghTiQEMS2u52zd0fG8JYkKT60unh8e6WLehzLw1DpMcGCSq8FzdOj26CUhDWQQ
wZQKXSjrXEEckswKua/lW3TjdgfomyVsNU60fH2VahXiNTit2rmGwZZAFdrSy/taNHPJRdOh5wCZ
9kUEtVaeA0JILJ1yABILgmHL/cIzYYNIt7xE/MFDypmFso7pL88D8gBwCy3dLCN6YOblmzcFui97
gjvg4Nq57tL3RbIyM9cXbMsRnCZHzFDOvObXKtqgcT0NdqocjqDe8UbBDTDXnoAeyZ19AhfGwPVR
c+wVUCH7veH7ip3QGmUxdhcq+HaAheLfm/Yf3gEptnZKpd0OzCdzcsHRGyIBCj6ac/EOMTWr/ZAR
+4N1qenaLD4xf44MJX1ggFhKctwIqJyVUoGMkNAN/oo6o0DAEx0IOxhgF0eZ8i9oRTvsRN7ZldSk
BeMILEn+MvO0eb+Bb3MbZlqGNhQzU3/0JknpcZX79NrZwojJbfn3Qq9UW5txkCocA7jDxeUg11je
Cwx/mslCJHmOtXMJ1tWH7zYQLt+1OmdNTL2XGydDBNoOj2NApMVH0Sqvh+jHUZC49yGOjQWLv7cO
0y9Der1O5Awv0oB1KwGH+YAkrHq6rBrbHjkznAbONv2U+32sOvpuCn0fRacJcYXoL6p+HS5fcJRV
UEbdQwEJhq8N732OTVzlp/ygeijq6X4sFkXT/TKzkdKoQNagfP7VKIKqgbLjCDmfedlb9v5V5/CA
dkiy/lS33EzD3WAMmQvx7vUocmF9B4xGSeA6ojiP48lVY55RfwEdCNxblW3vPo/aCxElbZvd0Tys
5SS3AvyFTLUOGaRzPsQAVrnP1k7F/HhXWz4+j6Xx5I17TKZ2H7i6DhZZ12KtyrlGiPv9CuVkzaKv
fCJkrvnBJiQY6/U1grsYnAoAOW7XykmmhFQ3V41TqhFQWB1GRpgve2eMDtBlfaYv1vKtUehxq712
+wDNJ4cYjqs54dteWV/NwvCs9LTJD93V2YmjiaZ3bnUDKhbGhwBn7CnFOz6Fg0L9ubYzxLTNAG3U
vBZ8i4AnmtMj4I+n1no6Gw+X10GHrnwNnqZC28Cy27LrY9uAVV8/LppXxUbpVFeShSbMzT10IZ3o
Yr17RgWGj3yffYL2Iqa1kQr1ELd6NQLCpsLpr4ZJOinJb6WzNbo4pVZJnL4f23p0oey8LLcHhNMJ
TkxkQTJx7foVhULjMbDsDwp6QUpqIKdjFBE6+SIvnx0I6BEWprMzhDNu2/0iIAvTGfRTn1psNpzH
o5jznlYel+s4PPQPqDNL9H9qDOJ8EOQEm9lTx01y8i2q4KMcMqcFgmTllDQdFhz31dBhJRBCd16s
5PUTYefogofFOC1wXYz6K+mDc6RQxNHwJufwjHMemdSBf0o6BvXmaCbHoh9IFEaNAriXxvs1kRFX
CfH5cV6oqkNOo4Mu/Bi/fY+8p3P0L0kZ4QZ5VyrLzZZgFzbTDxLJe1b20VtNXyRCNl15sGwp9Cpi
oZgxXLU4xzd+p9ccLS7QEkdcn41xkDcOk1UA9WRxw2UvcWsxxfyOuRrOra01IYakZbAn1xUsfJVO
l/d+vudZjfWsZ5Qe7Nb3ocVjiZlJsuCe+GbuFqALxcjZwp2Ud/QvohwmF9rHP/RJmcNDVvMDt37c
DKdeTdcFQM/g/z4Yi2Stro11sbPb2XVqydeN0AXJdl42WH3ZScOlqYYVK+Cclz5iilzeD908FIMs
ugjR/DguJw91BZY6xlwPMRP7eQDPKYYLD4FBnwq995626ir8VMsRPscIDxawnfPcZOw3CMIbj3Ra
Jh75SnXwllSCJrETpmEWwU+dq2ysZcNY7OL1/+qXGjcmMwpvU+P4HaMU4XFDGjPnJYivd5YcNHOy
lORO/L3YigRQ7jqbOD0xl+u8/8QnUt4i7a0KMuLCuYJRS7R7TSSj4QSB6hRTn++3yc4MIAtjIQfM
UgmQDjhRXv1bsYj3y+poZDPM9EfvvvPMYf0HuSPHE3/twlRGF1C6c1y9eetVQyGB7Ipat/qeavK3
90UrKpOFmoz7wSv/kER96a2jIF3DE9Z7CK1jN9jQcKAI+69trsMi0pZZ+ccrP7+Az3nb4PWeXXRR
cwJU//caxTtxOTmaM0lmbjbom3+xku3sXCZuqRQCid5I4fAk1fRinai/MjOALv70hDT2OXurjPLj
P+B2g15v+GeyoTnzsfCKCmSDvf4AzzPYv9vkRpmdf1DkwtShkMecRU2IIhVzMZzj1ZdC7jhXuNxg
L3tp9uA+QOp9uE0NElGoeKcx44flZ2qZtWoXvlf0qBhr65DPTAJNz6PsKPoI3V//SHJCHXrz+i6p
/05ipmG5bMkL71Pxg83FNgJpix2jSFH8S4aLo3iR4Ak5ekMsB4LwbL1zRdXnD6Bb5rRVIpnvhKKl
jADB/jlRp39I2U7fSAihhnkl22QcE5BfP4vKtORWzkLzBDsxU35jj3adPTVO9/hwfW/2c4pzg8MY
wddATP/OqxMpCEMuX9cDwlscPFrA/YhO910NCwQXHKsJihNVePStsn70a3GKIidOQ9IDhRu9yoLU
qSMiT+aTL8x1jRxIapPDEL7Bg95mqkItnsa8BGvYoc2PjnATiVgtoEBUlkDdZ8aiO5vL6HGbQsEF
+iqEZ+iD3tNmTPJSU8lpt9gysEVNng/aYQHjaAxUSte1WE73tZ0hi+1oXb7HoT0zf6xvjI1XWnkc
6t0JlgdbOdskWVXfbOeg6x8Yntg9GRWNNPBWPBcDw7b5aTVW4h8eJwk//l/nn2oodZ8kIEYKWsaZ
cl2P3edtRvCUD43aI/OCB5Sr509W9kspRgfYnRYOqvvqoCX0BxA2pUqm0Phir8y3heON03XvuM/L
nhz65eQgi4ubHm8sinpmF8IxLr2bU0qZjQWUk2r+cVQU5+O4d1cUiCKeAgeca4M5ccb8jvc4b1at
xu/u7SiiTsjZjtWC/Jr8UXdZxzODZ3b4QyRoIJ+KTtSF38f++lxqfB+GZlUY/Plg/6sY6BRYi4P0
EsnGjI3x43swin4G6LaT6Aqn03bVawW6KUPrYtvBTPRr8HPM9tRPgIMFfpog6J5ePtGQTkybvgrd
7JIVpp+tAiMBBSh2aLq7R5BxbNJibNw/5zaM+Ls5BbNSqtb1aHIjF0NGcBpkyboEYoEkwWVW1vZ4
o/vIRinehA0VymwJt0+JRuKIDfiP0SJXAV20E790HuCOKoqqwABPSpUNtuAetakmDi4qphOi7y3Y
8cdCV7wvt6FnLF4sZZs0B3XdLqlYnLZnOFhilPSXZ2D5DXEeMDZJGhuPBR44XWug2+T2zpAlQQ8G
/i+i5hCxf9n63z+Z+ULqaHVb17lhomxHygKaM4XuA1aJX3/gs4nGWIS5QrNyrIgVDixwAmgojuC1
AXMPJ/Hu8uf6WVfkjaCnCyAGRTbaTxF1uUyDR9Kf763glEwxXJ2zaxON5mE8biiXo5MobNQhIRMf
4U/+u4cYfTUKlCmQi0G+lz3po6UBbppHlTPtA3fo16qczjUBtgE6n41EP1+BsiCSzRnOJjfYyk29
Ojg9GTR3+QJvTrDhcXpf97I7HtRmPcxqj0K994tXHnNt/0zA1tVm+2P//efDb9xbruydNFzakVXU
6KwaBVX8jXGmaafzwscKv4Yc5l84mXCMTyh15+S8DQFmHz2h1yTE5SEXajCQ+IAfqxH+Q0/P+foQ
LkYxESaL3NaSIU7M/cOQ+4VKbbCYnKu3Ym1SVoIV60Flxnap4IHuc/CgiRkqlJhMslO9RBOTmFJj
wltmot9wiDE3FdunMBHOXW/RuSKXukIdDXoDzAjBLkJwwYZ39BYnHY75fqo0407Fuq/QreiIPK+U
ylE4y57JvBbAmuvjdQk3HmL5KleSD0IgI0Lf3YXabFd7r4E4MqQkCwKKG7lQF5hIUFMILMmc8bng
GfETCxhg4F4M5GAH3Y85TcIHAzC7kH97XnQESAe6Pm9IIvZNg5Sse7DoI+oBhg5r4chMjI7c4nHQ
IhyeBTQkrDkoq/FUFlXBdACBIs3cd7g59bskICAdfgPnclqUKkTP1aUBco5cqFMHFdJGdS0yJwPh
NEQPQXbwEasBt/wwSRnt++CyXSWkdDgxIgvgucYdtQjzAJnzo9tC2SZls60m9nj4YA+wr7MekCd6
Khw9cRhekSIFfv0rzJfOp5AKDDI00kKSFVzR3lJmLZqUUqx7ov9dTJ9k77m5b8lc/1EOBx9ATXsh
HwAm6tbbWRdV+ayvEa/PkHzKiWqk/vSKokugsLub25fonwyXAakGB6QkpLGJjzqbJBysiF76hZoL
qADc/+TtETbq7wbk9SE7G9GCi0HaneoqNzNwKTMKDXchI5EiKOYpPmq+yQAhNUtRSQw9RL2A7aWh
BSyUwpGC3OlDZ6PWgbGn9sTm+NhBNO3PwbnYUvmuSsu136LaWT2dOGToHOMgfrlyo7dYz9yFLFDc
CExDUy3cN7OT4E+3w/oawW1/6/188JxKFwdXvSifsz93piZeZOsGgLrrBlqmQWRTgE5BwQe0dNvF
PefdP1SM0t3n4bJdNTfia2vIvc5zikCu2pemKYbq6GPjl7l3NdliJhCCZLxVNBH4eTaUVLawc0pz
OD3KtD2Kbc+IUEaRX8t8TN8Wk/naNRE9evYUoi4F6H9eMDUI41evJlLlttgmp0tQvtrMfeg3dBO9
srQrW0faJxVmb0fUA6RK/5H2611HCXPTo5DTlFLSW1GjU5MNvMRKajS0ILaHgCZnPcZADzPU6zHk
JCTwmdnwxzyG9+1WymlH2+Gs4O3lg0cHsaLOM4XircFtUFYjxVkbIyzHsmmdo+u5gkJDT5vzxmJm
88NuSRJgJ1Vbx2QVSWIEaLQNl5OMHBj6K0omRZah6c0BK2I9WjvJkm3XaOCAPlBDxp1+FK4JsPoS
/vbU0MTLUhENnYx/Q0Tw6qWmm2Rz0OYrQ4AruiJlDfQRc/9RkAIwzTCZIO/kgz6aJ8tdGF51FRWU
l32OXTllA6AvloybgeFvMiW08eegWh0R6exJ9yCr4N5IjLeu0EI6B5F700CjmBX9ScjlGHSh7S6m
Y8x6Ai1NgVrG+2A5SxHIVYzkhLs2m9veIjOJoU9WBAb+HZXDOzCtVvaz+ZpfA/MjU15zRcxaI+uq
qKuZnJ2BlZNROVHGpVodwR6+2ttJPpMzLTGvUeJ7s66M0ZfwJ4ikkMiuzpldJM0/Fe0UF91tTPAt
jsJZwVCfGoimg+S2z80wrXoxjBLk0fRBJI5oSaxC+OWmlKtv/4ZSFShbdVCbqtsWNSKXKxxwiXxj
bjAD+ZVs8HU55zD2mqnC8YhFdYFy/quRjwDSI+NC665JhodXNsRl4KjnKN6AtOye+rRXgxw+5ZU2
3W6d1MVD8jouGBTD4WAdssMhliqnC6gt1heDt09WmbwqxWjcJEQF++WlmTmH6gDFIC8AQXsdDmPZ
cIZ6H5jLFLjh/gyhn1IsfL9VDlxZm18P+bCKSz64mdvg+XbWrCAi1wqgNmNcuqv/RVdT8JHoOdna
g+E4/n4/9pzH7xGwALx3L06CxZbEA2ffOcBN6ckst2ErdUaLQrZyiTMqUp8ZpS9yHq7Tpm6ANoCx
4HKufn0ftrIA35z0h/R5WVG+XCXsXdhJsA/lrr1BXtVP1MFz0F8+i6YwP7o8phCF+gNSrb0H8lFR
G1PNTm2ZS9AlMsLPNsjjY0AXKcZc0p8gaBmfsN7T4JrLjmD286SM4zr3gOYrapb4vtoyhdeLHpH/
LtEtFxS/RvQpcG5UBa0PtIsd0aieFgYopytnouLLhvscqYve+lpYjTKVXPqNqzep4J3HKbvRxYoj
+2V+7xG760gYkSUt0fhJ0ubCVU4s8mpFvsZhD7cokfKFfbkO4wB7Zas4zkKwlpkuUYvMTSQ2DWgz
im+cZfNJckqV+dNoN8MjHlSeoIrzk4O0l82K3hP6AOYWx3Nb2HEX9Gxz+i6y3G7GuoQewWBn8lbQ
2r9/yfFqGpJuaCxnzS3my1XUDEHbRfT/rGoWsaDDYif4Bcax2BWTk4Qf66D6B4noX4dP2/NIFJc+
4AiO5I+toqDN3V5tWHAtfnJ/GLspO0OZB7+ggadu38kkfeER3OZzx75AW85G/dH8LXGO/CuFrBw7
GUtrQfY95Rh54LZLTzvrIDC+fuPuknqLNQbjdpUcQVn3cAttzZ/5KhZ2CHqzENBBHCtOYrgrERcO
iR1x3/KqDVQEEu+hYZ/995yEQGwH0n1ft2f38M8W3FH2Ac5UDOFvF2+7CRL3hw44W7GZAjsVk7Xn
AuaVDArQ7GKsarFPbLRoWxm+vdAXC+FxB7AvV3if1DaQ2YoOf/R5nTZI/uxsA2f3dtYgKN/Mgjpo
fGWgrZBPoAXhNvtTiMsvlDaEgndKS7Qy+yfyEMXyg55/wBlDk3JmpkUwQHZMVQqu4emDWy1p6Ry/
+x2M/jribeOBvnS1AiN/u/VeCKaLB4bxUR0B53MDYd9BhZCIEffwC0sGHcB4SOSUzsAIJ9lcb3PG
foJ14RtTxlv52q+8ZUqiyj6biYOkL34NQY1M0agsMizY+tLD1uv383OLy0mB9ATzDIhi4paU6j7A
SNhOzUZbHYglswaid4A/faeIXwTez1Pxe3b2vwQkBkqd4QcVdQx+H96Xm7X4XAWihcrVIuUoU2VD
P8hrmkWWqdO3Km8GYNUfLMGZmq9LjC8UZu5YGNxKh3sA9u1qI1MTjTE9XT+zilGqXISVnkETXvUd
AZLaIiwNTmEApOCcYdh5yfCKg8HNZ4wKH0sNXz31xgINJyZeiAbO/8mPOiLjv1qQ9CyxzIo1yPAr
T6PL65T971M7LMPZDg/CG7dQzPZ7xoei7GBsHe2mldY+uY5Ktxb/RK2Z4Yenx5KAgux03r2pKsTW
suEKeXgwdN+yUN2zdj2a9JIpCiCKpZd7H5aEiN72sQ1XZL1HJm1NUliUyR9GpuxKOX80/1CiN+a9
LS19UIEiy9+6ErA9gynMBgJfWTnHn5ks8uxepWRoG5OtJjhmUqRnANwHSle/yUXPmQC3aLG2onIv
XtSpZmP3v4ElH+lpFyzEye1f8eJrSsyIlNV3VNVnujigdmL/PU1Q0JXqBW5MIdxLnppxlHtCHsG2
m10lgz5T31HC0WDAYkBa61tfZkNJMj7e78l8oKIVv8UwmdEqFuGSbPQ+y7gsMeQENyAN0fOTAXdf
+RI0kufldzQhMzel0OaPlXI9YjxmPr0dtELB/g8GQEa4ZQ+sBi+ojPfGItzYlPQkjCJJT5rFBvh1
bxF22x+KcpHIZo7HTZQ2mYLrEKDd1+Q1UrL4mPnjZ6P3KPYyk4e62MeSv5bDXmSIVkhYM8MrqXRH
8hbjnaKm1cAZP1NFHmtRt9OdSEDn98GlrnBGwcqg9+fjpSWDPP3iviG9mrp/p1RYG/Ot5YX4W2g1
H5xT3kwzw85ZwojAWWxQMQGOlkJdFikbED67xjlbGUwtF6YzTLRAXu08FPzbOCeX1RbN3BQHywcD
KzQfr+FeOPWhZo/B4F/4TygQiL3H3NyAEA8JHMTsmMHurSTszZaUKZw4nBlUHeWJHlok2w1WlOju
bSYm9/srYR+iN3gpyPDU9U0cXuSMiTWZswxn8zqt44b47y3n2JaCLPJZWaNVQZoaeBLhDNHxPo2I
CZrys5lEe9La6L3nfsDWntqNioT8bYfwhQR9YuTYo1Ste0ZKHzspdbaTSc3/hmtujMpnXue2m4PC
54FtRuiXm7AItHvwbKvFq4/DtH2VcXZJz0cPhrtXj8c1H9mAUWdteCVZD8PHO0RSQrxzLY0DButH
Xl/jSn3qTSTjhch9Mb4FXWb+Ax4kQiEMfFeAg6gRd+dJ+Zzba6PD1RLNEedVazy3xeEGVHdYCh/u
sUdnw+qW+7TOOPf6nw+rGSjnpIsB/ZxtwM5yNZgGm2/JB95HTudhtHVNhA9bDX9GPuw0FzAytWvV
U6acUNgiI82ZYjeTYZJtuMfI4GFj7a1JV3U94iM6kfQePCZqx3KR7VmGonG3zGaf8dgNKOCXfpba
zS+n7yX5/dUuzXA0hQc7VlZ1xPNKBpPjZkEpPbpNvEnr8z7T5j/aqZmQ16wUJS8lcv2eKv2u8kQN
3mdprorgchgkxFHFF9fHF5/vZ1seY5qBiDqom2pTmfWFSb8Rf5hMA/QLC247x1VKFqoXcV++5ro1
0OXakcVy/JtJBLoanql/9dukrHUPbuACjlabVNZyQ+A8v6ShWb32cpr1pHCWYzqGtidvZ00WYFWI
Q/TyRJLUfpOlaicA2i3NcN5UtOIvYx2gANksO1y0YAEOGLPuwTk7Q7jkE2NhnVJpcdny46uP8tCH
wfmU1w0dt6Nu5xw1tBQ2Dis+PM6oo8nXZ0yWdjXZEPUAqRQdR/yJd38K5TIwDO7mH84zVM/PSGxi
lyRDduONMLgM/h/NHUVgWWr4V4tI2bShXr10VSdsyVcBQHKjuUHjwejdf5pjjDrx9miAKGo0P925
9jVXSB9XISsjd/6M+W5k9rCFpHIMO4bwNsWjgCMzKvTGOcjtG5ysTaWO0IQ1BuwZdSMu533/O/7w
cbXD3GGeuHy5yuvubuDCVHFktrdvr2FA53enydOvDrGvLMsmMp//uKFVnY4wICpWi/OEP/IOJfWa
5EebcAhyx4WO8CiV0KrsSfaH+gsiQ/FyrcvB7teqkdGvb7P6GyEtC/e8hyvKuurhZvI0hmLQI3HM
KagcKLemVMIkdUHG4qV4eg6jcIn0U3aHtziRY+wLj49SeCFsPN7KYXQfLbK8n36UvOh5dfUMlXdf
md+iw4i1pJB92GMancScOOQs9jYVgfu8cNoX8lRp5odK2iKR56EqloB/IAPYOz2ahm+odiF52xgN
HP2XCpKDFlW1NGwWaF8vpscppjgBAuDcCOYbhFoSV9b/H3510UFQfkQmWuGsttgdsgWZ1s6nFHUB
v+K+K7f1c3+0s2KwgNlHsBVNftuaout99LJEfPdOzL2TNA0KKDWQ1yXJ8OXctNujnSgl2e4PQrK5
Lc/o7sM76Woq0NEbjn+3sDXIr4KTELYYbATvgSW+tTqFULZsuQpSuHBIfs9ihi+J2uJDhiYnDgEZ
HsR+NjS/a6gAphXaNIfajdsUKSZ79D3IlP4DZn4PWtg+prwPVuJ9c3/kJxd9ZxTx3M6GIfR0jIOc
AgE/iQv8KlIGdvnuwDfCYoODQXHb4T9prpkiLj49tOyqe+KuEjsVW6e6okr33ykFgKqSiQWwXDbZ
r3QcfGb7vMAvBv9LadCo2EzAOGVTWm4UCwHn8+Q3eMkSeYjq2+wa9XLjjUffTP8UPj8RZYbPJXU4
rNqm+CuN8QC3RvAZ2F3N6qRlR7lwezIZTb1PCCwhvygJBmZuXXIT3D9iwqLsjPDdJChNrcjCXPOq
08Dcb4FArS7RXK6HoNteeDLPtf/jC1d2jTO86Y/NcQGxPMVtp4Cd8ikrMyi7bHKdOkyPxrY7e/Y6
JBllTTHfVNHjMXun0NHsRserx3m9mt49NHL/2CIWoRTxbBeBZ3yHbDKaFu/9bIcfWEwXCoob4fgq
03Er9ZRR73/rfWxoEcBWViFsmhz6sVChtRJpY2u+OvCt3uHmLIPmZe7OhIOssOy4EufKMylzJoFq
wlGUtuhXIr8o42TM9ykMED9zzwg6qMLHtecQhCUNDdv/lLUszWjSpMAtc+zGzRgWE6bhwCeo7nh+
GuHXVlkauWqdLgZnAuHhGiEsiHUiRsqt5FTOSEuOi51n/8zrXFausOlN/7XTHBrIkO/t4gpXtEmH
qv8H61ta9E8NuBaOABPvxq/+jiO3RRo+LSYYObGPf0DNiOGriefOfoK8rkDxxuT2wzktHlf2FV5o
dUBaqm6kFQEpgl+HZ+Cc1+Ny9JVIxzTEw4GPG9tI+8tIrGeGauJs/RAvcnPekRbExDQ/gw5WTLXL
CDaNFW9VK+X2egc0LOb+4LDaw4Xfr2Q/0Mk4Aw+EqJ8xDzYB8SLSSYBpDHC8HG86zWz+4kh5U/L7
gvqEpHVa6wle1O72q7uJa/T1tVE1irKd643csK6F2aVMaOiUo/neqezMzjadl7ee9/Jtk2l+2FR9
5hmOepEc9dC4eMwZLUgBQPpsqqut17OoxrCa1LJ0CKWzZ55Y3rcY5OKm9NIGs16O59xJYU4gY67F
1wGuMh9Gz63D8KsUI6PiIhTH9vaWiSlgfXoBmyW/ZZo030saXD2M+C2Z95Dz1oc4GU+GMwzpQ3Ea
hirJ2VTfzoSBVxewprJduqGd1dwyVK9/Dk6fGbyQm7H1cS1K9218dq0jSJbkCBJUhEnqvkSl1oUN
4SrE9H3YGVz58c+VNGHuc8x/9e1IOET/m8+Dx5HYUQh0/q5vceWwyFSr0RPilSC0z2n2xbbW48Ul
DDYsvkDuB340XtvZ1rmHGenAXg10Lf6cQsVLCY241oCFbWf4MQ+DAhz+9YVFHKbN3I2qDDi8zcdl
32chGoqRRsnLoSTa29fcSVLlMZj3JyVGFzjvHO4FXVIW7qeaDdeVAzPZEjWPAWbwPCJtnKzg9iPc
CkHCh3h8TajcdSoAln7CFfCiGoB5Mp7q2YptKmE/e/uxn+VWLmjKV5H8jVJeAqXftRJjdDTejki6
LUMGgBae5ntX/wqdfXe60xgGg+c7zApNgOgOxnFKtOVZLN/+bnTabTZGplxEjAD+CBlLy5ndu8vZ
MUsvVOrXQR1j4xImoLlA2AChqxiYAbbUhuLPOK1G1w557UD5OScdxzs9RDIKBQ9ArRsawBDGqI2l
SGZCMy/gzF0iSwFRNi1SF0KS8i1WaSA6Xp9bTsJV3ZeB5Laj3ckrMfOOzF4ttq2EyvQPUgaqXCNE
8AOYi9O75VXyl4Bcka2MKPdhTVJJ1VnQMwRTtZLRPVisAPTve4SkAUEmbYaMiR5AskgFyMYtyzpu
oIuU7YBX8Pkifd8gQ8fHvUD+C5S+fMV56t31/F4p9yeHr0JX+iMVOSESli6NSFUZCnhaPi68Zniz
rs/g7GVBc5CUpLDvKO0naFm3dzZjLEoWcLYV18TpLk9psS0GpGK8EBiM45lVkbQiGcbRADDJGYFD
bxiheX1kR8GxvwOOdZJ6LUDr2vB8i7U0FxHyIPcTAsisTYJxnphWCp955hcEvYppxENJ7CYinU9j
IvwS7RReGYt8VmfIdmCHUqNj9/Jf9eyndQZWibIA3wpDF/2L64h9k2eB6tra9m4UORTRMFZKzC2V
V6UGkQEjDbZmVHj5DcRYgdAZ6ntnLwVMjQFr+dKsJSXWKmEBzimrI776Ay55BXRrvG+1bnSA7fF7
LbN83PFbSqgor7xAzgwgnrFU2P2d9OYZyesQHnX2cjJIR0VHFyjx4xfDqu4kJxJ0yc/kxHlwGuOL
BB2LFiGwPemOU1O3qOwen/wOJnkm+qooF0gqIlhxAdLG0kwe4hxaJLOwWj9qRBdztR+asCyw5eDW
rTHouPWg0JGUa1AxzMCVjoMmg42YJ1J0amjoZFSGDE208s6U+XiUeGL+gNq8PNBHSm+fJ2uAWh+x
CKfGFedmL3KKCU6Yg6znxhyjH4s7JamsMhTzBku+Pl4Vq+gckLIAXK84qO4TsOY1ifSpYXmmS1q/
twr4fldXogFMbvvYmHT6rtPfsg0NBbBHF7S6rXxFx7/yHplt6YitImdpFMeMN9AjmNKCx9Iz+thM
1eWOMVHrE8NpLy8G6UjKEm4dQwrEQ4KXLIkgwlVB1SG8JfUmaAjcC0hHMMOKo8fyMVHUga6f5BVU
6/oEQcPzESI5jPmSAzDAbm/B+U+4vdxqO5jX5V+pOtCkwH2VPiLsXrGkSgRH6yLKeZTrWHbxBJsy
RFZuoVICUw1v/t39imuiVddhMhas0E7S5dn+yWCkAnYd3SbZ6Ufylh7deZ5ZmwyuaYtn97BRTl4K
KHNnn7HtksFBgWs5GUpYTaH+g2HQtpe7+Z66UcPDS/VJn2ttqZaEb80zprNhXmCoc2lCd15v6Mby
Xhs+Xv8gkotii2iW4vvPlGeCxGN1clV5FV55VrdJQRPBk5vb9BMILzjkGdAoJ7ehJfrTYrEl+e1A
XUR2bmrT96NKxVeNzSMr31uPxEdcj1uzrZVvqPzre4XS1nKdc88+FmCR7tOLXQmveIiWz3korr2y
9XnGLl+L3QOiWjQ7Rd2aofdK7t73o9/vzFbN7XYbMIbSal3wOd4p71B5PATyn/CbSJsOn3gcpYeX
LjyoU47XjyBk+qZBvzJ0dUgHUAVyQCxF8kkqFV9oCxj4pqBaueysvkx0/OAp3j9kJdV4hJb/+VS0
mEkKkGl5ib9qIsC6vuzNw8RSAcvzYJDOKaKFbco1uhrzX/Ufg21UJmluQmwZP+991aQdBnCP0TFJ
ACnBPVT3O4wcPymg+rv7E/93Hv/NupH0vdZaay+9vrSYRe1kXQ4X9Qi9eOQuylZN0rawiuEg4V8F
/tfIKuMoXNfs9fMi1EhWHUpv+3da9BuPbb2bu9EVGmaCk9CND/7reSQ0iyi6YDtwupvDwVQMovcq
BO3khYBkWIWWM5DoxUdlzCXL5ul3VRo9DU0rdj7FZ1oE8wd05EGD5xGWpARJwNzlZKcd2C90CB7O
L5XfeuZYzdXvtk2VBZFrZGiAVlPeeE2hlDoYresLSgMHX3QAaxLg3NHAfKhp3qJ4Fpe5tUWESVA7
O4eekgM4FSk8XW2njvkr0bPEC07Rbi8xAyoZkr8Ujzr7yT+DfhDyd9sVpUmeZCHrNmTLnAhuaJUd
3Q9kqmNAYRqFdrjSlpZqe67umBLhye0EWs9/mG6uY7Q4l/8DAhjsepN1d2B1q6dPD8sdti9jfKSn
nRGLGi9d3+/29pBBBsyOrUMj2XRoz1FQOdbxT8RcGmqY4mSROBOO9itJzgs439CxBtA7vlvD/7sb
B6aLq/6FmNbEfrkfGuz7e0gfnA9AMOA/IbT3nk2IYCGCiDyYJb8oDi7V2xV5xMl0B26654aVqCMq
O0JyBrEFvibVuhoFAGHbs/cZ5OcSyNKZRRry0AsRh81oCgLV+jpyW/g0NRbeeIxGZNRYZINap2Cc
rgIKeM2tnen/uDRJPPfbUxaxdsEf1aIaFLMqzsOdiENJOS9ZgS9Y9XBHsIpz5Q3zCmjKt7SRaZVE
g/kn2VPPgnQEgVoVjMfMxowUz3Y36ho/yLWssnjfbApgFKN4Mh96GnOwkOo0dww9xpxyjrTZUwZO
K4sQhWBeLCgJ0FFPAJHRWidRWkPHnMdt1DhB6uBOKmL52GvCUPoJOtksk39CksVHRg3NjJ9gY86p
3PNOc6EUM1qZEt/QbZJZdHH19/FY8DMdljuWAi15AS4PyZQFIbIp0fxtksGjKA9+ItArlZSdqCb7
X9x/waT5mjyqS8iB++i4/cSbYEylr7O7AYGVDCmeXbBrUCHP6sWlNrfO53Va1c2O8wbsiERCrDgN
dAFVd2toocXWlhzXPKykw5FCIRDx/EmfMBchQwJMRGG5N1IE26xWloVrhzmbr7IpFVaebwmeiGhA
5vhLS4z+z9Vt3+ozydxSJDsSFfiV3LIU/RRBL4u56MGWj+E1shVf24SVCOjeCU8GfUQp2MKdj6M7
WW/d6LVR2XuM97sAl8Q+3EHnziHyK7ME9BSAjhSrRTx7Z5ub0AuTV5yjw0MRpnTixYT5AzdkB+Ih
AEL4tBHjcZ7T40T9uPLVfj45hYd6ssG6+uKofNkdeCCAA6Ng1B9gcZb/1bEmmqPXFsatOOhy9IW+
tQ/IF4jxMnwdsSqZqS1vCeCvtv6fXrMkVTliroS0QlRFjBxx/KKXMl1TjSRSOzw5OgaP33DnUEQ+
jtuWO7k5q7KsnaAMPlesGDh5VihgtOl786fsbE46Hedtmva3OeEGdHkx2cnsx7dB+GlkL2YrETwt
wfN6BRQAuakvsfJOkk9iO8pCAH1r0k3HePX3Wj5rNLoViXvnNhnNd1QXjiY7xSEX7Ewrw5JN8w11
5jxRzzmDOXtdZHabmHbHspqTP7W0iBrq8iPxRwrnJvkMrtkYjermWaTUE8idaXNOwQNBlVfKeq/N
AGXavhnfQ27n83OJEv4OULvVaDVy+NP4LU5V2n233XCnK8AnND5S0trxZQW3bPte9WCXkok29qGb
83O5AhAE+C5e/gWO/YV+9a4zfQikkjvLu63KapSGkdXoy/4XfLlX/f5U1CCpMXd8dHmrBq3ZPxpn
TVCEiAYAu8kwR1EBD6pNpDwE0Zlla0HAXO4B6B2bhfAZaF36Nv0scUcIJFuihCzk+WueSnwRCIeX
5zBxxAfsUpOvRy7ixcayV/82VBW6J4gnmLtlWJ/hkLUyYLNJZBB1A244zR6nKqAZmeQq7boNZ3vz
GmVrvOuLOp26DSHiDjzJDUYmVRa35oJRK5JHsIkPohVelJbEe9OQHYUa1XqIKrzAHm804PVDpHO2
iJTBgVF9EhJSri7qgj2Ilz+/mPmPjVN3aqd+zCjkKtB46GD1vZjRQCga0Ly4RM02OlEDoh+KXtMq
i6Y1HxA3qiF6Ia7P2tq9H1b0Q6rTKgcJYPCHdl5vx1nu9+wDfUwpkfWhhbpFDxjHAB3ZBVtRfuko
FqG92qPVMIIZgGkKTzWXaCkk6OMtN0f6R7KaxJUK+P9G6hADfHMfxRCmWIq3vDhtnX80Yj4zDSfH
MIOLKP+J5dykAKt7vq6HTBei7n4D2P4Ch0Ve0HhF0nFquFN5vUIA/OFXe0E6gXA7dRy4Ojf+L+Td
DoanRZ2SzDh9mIbLK8oZCvQP9bypuN1U9OT//UdnoOPjX4OzxIM8sqYxOJGkvgyi7cZjt1QJEtgg
zHUOHGTeE9AVjkwfgDCu7QM8jmfq4AaydtQm5ogpfDmPGNoT0AQ4WEkuntRGuJITn1ZUeewGmJe4
RnTpxPPIsUTAE3k1yyiEfS3bbTqiJeSXLO00D9RvvFqMOLYRHQtZjsK+Dgk5PahFF8m9VngFc4C8
E4I/BV+sM9fz55akYvFaNyZTXzFmK6PMRgsMzvrrnAbxoQWB5X0D3wVqcA7nkMnCiPtev8YRZcxj
2ohVQ+AUoW82faei7C7XmgRLdVaaSJCUzwX/N5WjxSm/zxRtUD9DnendWvqGApad5adeel4QdREf
Mvvkmms9l6OiiS0h8vMrmyziDBKeZiTxHlW4dlfsHqI3PcXynFf238mApLHIeh5m7iPD28Xguutw
Q8i3rNeSWYggW7xqGaD17g3RpGRoGR1N8DH0xz2TQ48I4IaVUzK0vij0rnRDKBuR9dj9pf31qDvY
jJbRd40NFlep+H9HgTf9Y/9uNRtk/CFh/GOJ+5bR5/KIP6UoHEm/svbxstKRDZMHKQCGp/y6v6LI
btndDxbRCf3TxgP9Q1BjPOM31qQKlFSwC4pFkn8NQ/cs4sI4GcZaCs0PB83cK6Z0KcHy8QS23a1D
4T2CUybr9Eiltu4xcp99I/fR2a/ubDpVmaLyq+zLgVQoMufpszVNju8m4S1QkljxYt5VsfvKY1Wo
a3OiT/V+XCnO/D4cwaV+I3RVA8x7BRUVehO6UqD/heZB1A+4325Txq4HBG2EPPNsSPS6dJCxKWVQ
xR7y1LZ7zKsI9Q4sDgIwcLBWfWvq49J1jqEjocE5A6g764w2pm2OehcUDzUsw98akzmEwb0qOgWy
hwg9XSVqyuW1+VQdDT5WjKROAQQm3R/boAQ/T4DANsyA7A85lEsrJfJO+zqYtk/rREuB6cZwWd48
V+R+frKRljquzh+p/Zqt5Pucvnrg456H0npCgb8Nk493DdNplvEpIq2SuEPNu1+7pamVmXLTtrwn
X1jWwnq+sXhcNIAoh0fnFdLflJ0Bkc1qWWe7sMqd4NrNSurNVafL3jQzzRFSvRxvhlD98QkjF4TJ
SAoYR7lxTm27hZzAB/ZvXY9GwrAZ/nefi2bZU8kwLHeCrSMYABp9iFOA21UkuilMBkVTyjCMZGz2
3LLyBvlczcKLbb4gIcylaSQdLpYdnkMCO8Un+gOby8qmJ9PwDNoPsLcrIT5k5e2Te0PA6PcL1J+H
m1g6XzgYRV0bQoGteME3AgzbGw/aDRMH7n6h/uRzGVxOMac7Wr7guE/y2+Y+uqZPNGE6kizNruXr
+TiCT+M95Bhw3GFDS1Ul8qFbp8P4+m8BCGzoccup7btaal/HIR4KKvwKWcO3xxzkza0QZWTBVRA7
tbzlk/aWQEBYeISjHawGZzh0wKz2v+64tmcfk+XKGg7s/imOa2Vfz/wjRHRbT+Ap40xbqLuK4LgX
vGr95HUZ5BRSKroQ1t4/YkhShQeIq5Uyq1CrCXhDT4TnCMvN/Ngy3HU3pyZolHwtpaVmoxcP3L9j
HhDSlGNOCJBoVXsEcnVVEhd5UkeDNfE1SPx3oZOAf2+vEorj4qHHPQ40MsIgKCLe2ZpOuF5u1Hib
P/iOL6DFwKd8jo3dGtZX2tqO/xshd3MbOcQ7KTr4wCXqae1r4v5rhiRdSW/vSS5B5m4k4bYua8lZ
w4QRsWKyFfnGiSc1FtVsQ7JU3equScohSwewOFKK+JqQsV7kD01zV4KsyJlPHjUK24FpoCjEx+y5
sqyiWMJ4j9YCqbG6b2mpHFPXNP4Z7WWM1VGNt0JWnZwOV/1Ou3XophpW+6a5GV80ogEcAnCbQEFg
FBiMqpRiilps09t++ey7HRge7f5jKbkpAW1Ygjj/n/8Jc1b5JdrWAdXMtqgImsXfIlhCeqrMOy+/
G6f9YeGM0oldiLjvlz96ESBR9WGHzpSNDtXsJgoLWiBMGpjlJdK4jc0x7Fx/q4D4fKfYclNcNXe4
j+ADOIPLzMN4+RxQan7ixieUQYnIrCJHR5ObCr8A5nBXRcbcyFmdUdpc/Joe3OupmLGOkURvyTAL
mIx/KrOwH1l8S+R/9uJCiFIfZ9aDvYeT7Fwc7PFG639zXepBZsOuRKzV+bnBRBhbyr7IpqUkD9C9
nbjQDWNbQt07GlOQMo0g14fO+n/Lbteq+4mU45+7Bjf2khaigdhT7GubnIMQP1gfHmeDX89tReix
atvG3TP92awj4b3PoV7QnQNc4tb6GsTvoiGm1RxIUwhcXY8A1j35WZa69SwHzCvgL2QPdjkli9PT
I8mKcSAlx4T/1Du8fS3aXm9p+qF92ZXA2ebF6PSp7ylc7t0LXIDrQbFtE97tv1fvmYHsEKSiaFWq
YWtUcbm/7aJW595Q17p7y1eKfC6PE7TziRZ2x/KYhU9h4ITWqHt1FVGTOrnifji+OoRyRlyN1UM1
f3CfMHP1xE4333Lz7AL3IVeKvPdopm0exGxtGAH7A3Vd+XOCnYIXZ1TpdszqPCaSstBfKxvrrKoc
sLDJAzUeXgVy2cdMLwMNnP5owrOZDt39yoY+4LhDVtjAhiuQR7zP+q/qCSXLSOekQLkfIAtMaA6o
S5DsYLkuOxQB7fcebCXCFoDJGeLXGruJqGriLBWYZtoAM2XwRmkBWl4xNMGjrgVwTsgGHNJQrdFx
FerYEImF/n8yVwW+464F/myfxRwlhkOMGeT9gHmoMyEf4mR5SD0ydrQd6KMGQdcETdur9BsP3g0u
gdtuSsXlG7NEbuZHXeFKG6spYbBaBjTath4e5EEZveW/V0G+WMQraIIQ6mGmsgR7vj3HqNGnzLZr
OmHfDFWMcMFDGOmyCSRZLzyoITBOJYEZ8kEG6nmteJfGGU/L3uA53Q48moNTBsc6rXxPu5iKi5Y6
zU/ncdZh2kMfeWz3a1zvV6h0b/zclexgQBQwID8ZPi6ZGXEN5G0bE9Mk5RIkapGn0ktcClYG06xo
MBVRc8MCu/KxTXZTa2o6mY5QjlNjzHtCxHyjXFQ+EY5quoVFtyUJGiuuLufkdRzg0M0pgwI+5ZXr
INOgMwG6C7BZ/kq/TiOeP0Mzoe5AlgS6N/nSY+Pji+AISckCNx2sF0LFa+1ibnvCPjSiX2b1mFwP
8zdU/Ilx64o7Qh5t+f2E33dmi5AfhfduC/VTLcuAkH3UVMNSmsJZO61fP4ThhJ3UVJasYZuey4qI
xOhXnTi0cxa8361eArjKSRIfOjeUamO6w9FdnAfE89KwfmBvWY0h/oRycx0uahcTzbcUzVWGz7kX
ZSEmwXVfu/aXr1Yf7AbPy7M21Pl1A5fq6oVTuKPR5fGn3NqdBHUj0EbtaDjA0FSJTVK3Hm1G8h6a
tqwBKksDhIng0UpkwLsmaCmFeinH/cpG8d9D1d7cTke0RaRRVU+HO8nsQ3zu0KOEua13UIo0inGm
qT/jB6SaIPWPPFBKwh+QR/0DZDwyVH0euEMgHNouW5eRAqbZEB1Z6Sujgkbg1zSn6dSMbmhDW1Ji
wEyWDmmlyPnpIMTudh1Y9DZblvBSseKDmG9mf7MA3vPAbXzhYE4Ck/7w9PP84Eq+hH7hoGHRJxmS
wqRx1OzQIHyXjMA2puD82/Kh5UuNQjtwy99KWBm7eVpkZz/FaaiDfVJE/LmRVlOhbXAdyDszTy9K
TnmUmgNBE9bLGR5HyRIcOBWEET9bCPxgDftH25WTjvMBX8+Q6kDfDLjfu6KfAtrvpXJzstUrP5AY
wFgLjQD/Q5++AkBZTUmNi3yKkQ3HQ03CYRofIKjdx/tlb6rj93IPGx+AIOMUmekG4p0NBBZzasUP
/zpQcOUYxV7ohbRatR6MAAS1mH/KWlpjoYmyT290KTkheHhUkoJVgNVHKCYeEP30YbbE9VdI3WZC
3XD1jLcN8c7GIk23w/uaZM+4UHm9/NaGdHwMIhimOGFaAwiK13VO2/s9WcE/BXubJjBIlRElr8ia
gAqubYvYrH5aLm9P8VL+++6AU0WHuku3bTMDJZRPD2MOi+jvD+8ZP/kBspme76jTxK5mRNpAuiES
5o3BCqvisI8BQNhG3R8XPkWsbxhspn1abVwEYIdAubnid6hYGlhwgLJP5iaOd9MeGlMWKxfBgoXE
1tiuhNBQkaz6eAY0NwOkrsdccY8rop4Ai7y3o34P1povkhI3plwyuXRvb5T7Kbzfl8g6FaCW1B5H
1gPN2MGcZVJddK1p+q7jvjbZrOAsutWAPJn0t24yGpf6ekUT+cKRM/wqYmHX0xx7Hj1TkLsck4YQ
f6omgFdu9HkPqzixW7Gn2++NJBnQUxDUvTPh9arhfl0mkJi6UR/QrhLv3ucdtDenwZF7sVZjwsE5
rm2BzwlQXhGXT3c9ARNHljYLAKEVb3DnBbx5LvltAtfJvfZqmuPLrTo1B4ZAwYtpqhAWes+bstCU
vY8FREx4fuaQdAMyYDJn8YV83zFz9vL8JNISdWNHm8IsvzF1xfoee53nULxd59UexFjbDE69y0e7
9AHjY2nXx2Y9j0GHW1lJ2nT0V0p5xTBzrmbFm655q794QX1Qy+7Rf/G+Zlzcw8S/gWt5SQRlNJR2
P5u6bGUuqqlwI63Rgf5/PJmvT+P+cy8Zk5PMo35HOi4DIBsDsBijrKMuNm0sIADUIGgAsM+3Lsgj
ekIP1TGgAmiBAHK8Jqki9tP+9aZjGnBzBJDAC0iVB8h/87O9+ZbXI1loQEKxSyj2v3FIQRBgZJBi
dd4Lx7vjabaorbHPknKYEOEUjsGnIfMizXSERU2sSYq/uoB2284hBNnXlcNNFY1Z1q/Nf0p2mTQt
puBocWfrUIkhDzFLB+tmPDXrkzyUxgsLIgrNwqLaClEwI6CpngpHbeTIneqWp4aoDrjv+Ky1wBz0
+p4HSNKAsDPcfdZqP+KoULoG5LRFvOz9XRdDId6lw0iF6QUtI6oCb8AGWrwMa0WsTDmddREZ3O2V
O9cUlqACjMYF9byPtZC20WMA0To2C0yxuaFoC7MIQpxRtXAIpeRiF7HAPFE9yXrY7EooxaSzmtwc
Bh9u9ceet2dTKEHpwjAnTtAzLz3dw02d3OAWgp+uzEowqIqeLgbvHuD32iesGX72L4ov5aptST+c
FS1MpLX4020kavHy/rJ6V/QXaZE84j0O1F/u6pl8vgio34nBZVbiUeYxWM+U+noAM2suoug1H4ww
JbSUWAZyOffKuS2cnvSQYpDOJKZLlkrCgdUaeY4KORDSt5ecZozyOmRfhM//rCmdzc1oogEK9Kzn
2BrwGPF/uS3IfeCc7sHjjmVQb9eJ4VoAoc7GycMtWkZoKueIBRHZSQq4rhQUJ5C+aiOAxWjzz3lR
RTHkC7Z6gbzL1gU6anqIeMQVGyQNyTTwNnpgj15lyRZRvNtENOZT6HJ6M6iwbb9eIPwZ2PpxP0jS
xP1dD6cnt6GdCEpOfSKMSIrA6PRRlzoOF4/EFlN39J+suPrUfxEpuxwhOxOd86LOwxlzRs19g46A
c/nlClsejs9NuELqr0p785nNlvYEEjpKAlNOn7xvYiPi6AWCQMmYOq/cWQQSfqJrt4wVQtVKq+Ak
w5lMO0dv+U81CFt4nkhgjsn2Yim6wlxYaqiItK2yd9RsmoleyllmrEdWkEOcp4ajDFO08aVLXhWt
akywpgK0GlhUPjWp6rteNtvTxTAAi9Rhc3j68lqcve40/p0xXouOJXI/xUsb5wg1YIaeRj/0ZcJ0
ADvaCyRHzvRUMP1q7FdguwJbJ26BczuOM1z+fvXOkyew4d4zFhgTWYKq4yzTCOUvEkAb7EpMp0y6
HhsT4lKk4RmmvcwVzIk+MArM+bujuZvGDL1TeSp9wYEozW1SpNWlCqRMCuum6W4yso4nhc9kDHUG
RvUEWtW/dnnVn39/CkaYIh4RcjJqxEBKOLRBGCJQeQin3iZIgWp3Ixp9t3PKoJ308dEyp42u7b54
IQYDTb1G+HpvMdTTQNw/j3di96+UrT5Rca+85nZmhxaFOUPhlZnPWUn2jyhta+udQsSH3ZFEz4nv
W/42MsnsxlajyoVkp2XDCASJ0LS+/M58kbp61wiQDpcfEn5Zy8NvWiirjV3UgF8ukiAFpt602i9r
akoFJtpIOjV7eFGgowzAsILBy2NdiOhKvtrmeEYrQeEgkthBdspR1YhLpQdxbXNn7IEr3V6l7ija
z/OOqqMuJ2OseIHKRWEy3u8v9cO4LYInweVwU+RcXEVl2Tkfj9nGJrTn5lARVbpt4rKSzCmaZM7p
SfOyT2XkSl4NsDDM08cHsYX3O9xvWdwJKrF20cuG8c0BYxPOsAkOXFw3988vgJkJG0BAcZDN1p3G
w4I8B0g8+zjlEa09cAejU/hkJTjPXr0A5GtDQtUtauSXM5YYO8PBNTU5SDVya1HqfLSrKKym0x8l
jg9wfa8dFVibUV1rACl2aFLNPlQ2u0CgflEiIUdEBXPd4A7dhxxo2IBjHkJZtgdSzIbf6aqYhk3p
kORFYwFWb/sxavcylLWNjmtKhxAm5ObBtr6fVKkYcIaCbdla3B7FFHL9wnucn+7TtjEKel9CYz4D
SSYFsCAlQ7LckwgiU0/tIzuSZDblUscs52+Bg069BBIhW+Sn4UfJ4mneEk1k0u8Ixx1PniEofBQO
wDR//lNi4M9FRQe6/mqBqxfK+i9j8Tln2QreoBfJluN/u3vBGvDUMuUOzCOHJGxp8JynzYIi3fgw
8zOrfXMm42CC2ah/vVNt/N/o2O9d/o9qPAC6Ieo6Zbtb+uil0+Nw3a6vKBftiyiQRtEc19Bw3SGD
ZviV+PBaS+MJ2i5wjIYWOoUmWhocUTR+OcS1dnMtIjBj/j03VvaTQyTpXc1O+4ychUsLXKNN+Htt
pA53VzPobPTbwyoOcjRLZeMVZ0oyfr0835wGXa7opKtv4BHMezMQj8p8uZgay11FGgWbikJZxMPY
9Yh+wjjb/ny4zfi6+eXREbsPASZecvOlVEromrpcVqPIvfwhIeYvxXuna8U9a4am22R3MpcwXl50
92LiqQngEglOhRsRGz4ucHeyyt7Zzy35dR4UbcCeiz1woViWRbq/+5SeRatjFQXj60UFukmL65QR
GIQUI+3RNZZsW8lwQkv4J1OwODlDPN1CfvjprjIPPYN6VWhCG9jrYrix/3Bjn+bljToIP2dMVjAC
K8NuOCOWxqXjgbYMy3urlVogA8yd9//fIGjKyuWmgiOJ8uPR8nkg4HhITqgeWtETlgdz7fFcZgI2
BwnP5G2zQnHDSq9/9qB04UkMKz5f6dOCVVO1k45dSLuqlR+wfPlKYhr/sP0BdGrl4AylcdkRixg0
W8TBXV63mtdDNgyOlctDMNj1duw0LpolpdGAVWmTLtFRpm00u9U/UQchLEr5UHcfbRRv2Tg47f3p
D/r7fTqSws/fgobwQiWWIqneSHddKZfh6PtYaI/eGT1HL8LWiH9MwVTP+sLeUY8A/m0Oag8tCoRL
7QmlT1NSrvpdtYMNMC1y0OX0ujc7+UUZSK50ozuOUy+2eYpxqMp+HcrinlgmcRPotjjEsWF8FVjU
zOhreuANHTnrDFuTy+ZoBeyOaa9STO4wt/B3x3rTggPz2801+5Cdm65jsp8OzwGe/VFwAbK7dEfd
T9EQFW0YR/EjYCFZhXcy50HDQlweEYDuWQBZ9VyU60YJ031sSAAqmoOXZyFsbjBmKalaFrnk7Ctk
mQitrKyateAOCZVR8C+u3lSHmSKY6/dgGVSRTT7FZq4F19HuAzTgEGF8GEieuJK2ui9bUxCC7ja5
/nWtCsw8pkdK8A0T0Om53y1BbkVSGiTJdMfGM1NhG9L/fRmnSfSctoe4sJTfIZHv7kv4hfmLCihf
5C9NdtxAe8dYEJ6P/XpJ+v1cWZMcSYY3AIgpV7w7gbZqW65wAA7hOMAcY6FIWo+9hNuAW+PZm4vt
BdTwswAw4LpG+KUumfIRhAoKBBT0U2R5oqo9BIM6nxzYmIxlCMCRMcNJx2tNBLB8ebLzhjpA0DZe
9SKztIEZZpcOrgBhiMyB37mj+tBD/wIaJznqD70bQJEBK5xIxawLvmkoeF5Pzbp932IfFALKd9I+
FZ65/kG8ecY3USu0eYo+oq0pDBugctz56dv6Pj59YxU0CHQt7ASyJy4A2yWyI5HGqzvJmzn3bk7a
2jyEwM5obcl44yBsGkkEC+4xkJ9ECPen1b70O0+6GD0v6e4HlmkildqboAzs+0cZvqBXEYAqgbZb
bOnjLH2Gu/zmawLL+A1e8bbC19kk3i5BlGrS9o0akth8xG0CxXhMHmW7o/plSsJvlWDqpSIYohjc
KcN0dAMHJRvNJL6K+rSj7/2zVbwSWckb5HXFN8RfpzCFSx+IVqileOWJdZGiBPISW0nsYKvtkNEi
frnB85JMVMvXj1QqbnCdJ4H2v7aQgmcCc6MyFUbSqzg/OkeG8erOjf25jBiFwZPx0JGXmIBoe1+H
fsJVnLjc1Pnvn659PaNyMBMp6fSWiClTHl/TySFXVdgzG6BZYpiWqi6lKGYtpcvkkSnrmdmOIn5Q
RjQOt3DV1yLOHu57/pQ+2P2nY/1tiR0UUQRD2HeNjdpsKED8WtuzZW7jxnB2A2zkKA4iSqNFYed+
6jjneKB3Qc1y0b1u69lyWmtoPBfrmb0Mp1F3IRLWCh3/1WPMWe6rmCRas0A3TW477QM1mdd29o92
lCsvrfPrtop1/N3fMR/6qL5Rnlt0dxS/uWNRmemLYS8L6+3atILaYhsW8jWBoTi2okn5y526a+3N
QnihJsRaOPR5VV+B+tVJEwIXpnk7iWC0R06A81HPiEsR5syrKRHp7RQJnzU5ZT7Gr0NaX4D3yxt8
XdOpqb0oisnDWXWJHwANUnRk3k4+VmrAgBj8RdaVf1zj5nheYQywYPRd+WcnE8jtFGcVEdtljR58
TMaLFGZZ4Gv51L+b98upSKXT8oegD7iYOEmjEsPiBQ4NdoTpC4xchqHe9iBN8DPmmGNJE8TzQCo0
H2IaBUYAx+EDG28GRQH36hAFykeCE8XTY0HuEoHzT5O7x8u0JMycs0shPXeri/dE+sDC4ZTb4X4u
X2VyUemIiZTi7MMXHCf02CCGbtTzq0ThWjK94VZDmaxwWk2Asfpg9nxwyKoh2p+kQS6d9WN5W0i9
aJ7OPTexngCI+VNTDAVE1/ttZ7+GCDGZPiGCcbyZnRB9avnGRLResk5CrA6/lzJzEJsylA4y3THp
du8KTLY4LnOJSi0FknqQ6IlPhnk822qj2aKlI1jJXxq+R6c7wl5cEBQcIm81tJrgAEosV5PzdtVC
iRMvX+l2EQdy2qAYro5JRty8ygTBgK99ZaHD3actQSiMgA3rIJehEllRP9/MQEPZaEQ5F3ZblzK4
O3/us0X1vZSholfVLOsUkRZQ7Dc1iKHx//Ru8w1DA/DEr5RjKzHXTNAH0CPU8+93ElhRRgTF4lJF
IL2MyAHX8XT9hhwOqzPM4Yi9pCWMbPFRp4YoK6pMyv6d7wVRQf0xctLbqQvCQsvzH84tryhOogTG
zgSU/Qk67rmbEROmPyporEofJlevt5vbwJUBa+Kvidyf8spTDL/Gg37Dd9nic8nIkPuuzMZGNC62
hB6Hf4nDIvSteUo4Ma9U6ibaYgQHihFHekrDUkyhhgvMfuaJpTu0viClKBhBPYY12arIGhT6Cb1u
QWpgaQ8eTjW0dmFIJEsYIoQdcMkT0Rd5oPE/9vGPbl8JczJBlHHMZkQBTtCTP6oVmwFjYO1EVtzQ
PDBbvTvjVJRrGHnh6OavK7ETj7f9dKjAgbYlXnjLjrQlu/HB2jm0H6QrMdmXVj5FZ5Yepp9AhM9d
yP2dkfEpXXHu89ML97EiNLguEG7PEMW/m0XIGvaiSrCt57jhsLtM3tAka8Y6xQgYaWoxoXQRqgqA
oWybWxh2zgqOJgMgAaBjp2k0BscXfmvuiMDZUmKqukqMxma59aERTnyf9Q+nhd0b2k5wxdmsBisQ
QleqRd90IugCNL6hac7GUo8PVZtyEDd3YKpyBMLudGCcp+XrJ/PzUBkdnQeVV3ef9O2Yl1etrBES
iynQ1ZBTNjgu84Pnet3OEVS9Tdxs9Wpgypm6ng+hrbq6WvUpSAJJXXzd6Xyd6B+c752jHh5hu9fd
B/OaC845xak6MLAi/PewEVdu+x7+LBt/YtMqGciN2DcOMO30msFbbxVgdnQVNEyQ26KAVuTXzpgi
oeI3XRdULRXm2Ut+1sdbG/2tn5jg0ksKGcvIk86EhKN0LUhNf/a35/DVNv8tHm6T3DaOCmeQ4ES7
tu/MpU8jRVO66mzJiM4ThpeORjjLa38/1ed07ir+kIYhqqZaZ2OPWpMPgul4ic3xlbjB3aRuf1TD
3BMFnbZRw1INgUeg/SAbvfJClpYsd1PQQDdraVJ7rbhqhaEeymIh4dxRl9Ml2zM3fhZsRjNd4Vgn
uMJEfHlzWRmxqgJx26siLYzAlNuDT8NpLROjWkihUt73lEI0Lwnhw/PAh0uO4EPyuiv9P61cIKeV
M4BmDMIhz6lHL6sFNke3mkHgNTEi5L1//vzXzgzx1Nqi2GtFe2B2WBvs68KH2Uk9UInyuLNZz7YZ
PfrhEyI8JmiXjSHmaZBDZF2IBOj2ZJtecs8WuFUlGCd3kIQTI8KqljY1WARaFBUtjsGlxquD8My+
ock2FmrU3/gy7EvxGdXZsNFYCLlPukyEYcHaxYewYZHo0qhRyOXiqfEMsDvX1bMfrDsHis6ew3xh
pZ7qQL7qWRzCBQawnSNTnfXx7cGNcF7n+JcSt62Wf+QnBduiGy+yM8XsL+pJtEZaiZXSoVN7El3y
6UfbFekSuipHjzkG/BrPAwCV1oOyGKZzmAmeTNkTuv/6b/Buxlqh2bc2PZv85rXfnnDGN0w+6LOe
Oh3hPXU+qvWY7VB24R+EN3NZ88Jc6MpLEcfFoHc0VNUo8kEJW8bnmwbJHWZmSbAeEKEoEK0rUe4t
Z9pS5gVDqawS6rzcfW3F9KcQSzKrPxTFsFeOQXFeHoK9OlKMUcU0jfb505wYkoWzZcub79JFyLeg
wIJJk/DSqYciKar2Yy9HNqzjJKn8cKZFlO2pARVFzjlCyJ6r/cTOpli+JvPpbnWfVhbesatDBytB
Yngd5uYAvQP6TwNryJDSc5S+tsCBOcN3liB4uZ2FEl9oADB/h8xJdM4u3Z5EZ1rHUn+k8yFyHgjO
3U6YhZOpoXk9+IYq63DHoUJ9W+0J4Hc7A/myuw9XtLdkWSvIGOxbfy25h0pcxYhWPQJiJxQuFBy4
fdx5I5AgzB9u82tSg4HsRBRdBGAB88EgFAZNXZ76/RxDRK3CJYTBJ2+y7heQ5ow5pRzgY7FmnQo3
/k1He7rMwLAUlLLjjVY/xXuvlUb9yJhtnZGRRK1oEfJ8kwJjNwY69U6Y1+PnwapLeM7BI7Oj3SAA
xolagcVSNhzHiAgjXiOk5FVEwndKbAH1WaqZ2VqkwP5VZfelNleguuoRoBf8JMv3zVqGzG1lnZBa
Y8VRdyBqQ+lGIZH7twdYnfDLGKoFlqLQ6j+ry4ZM7QjDQQmWVFn6tkVT7HWqC/dEpwnFaDesNQ5y
ntkH+pg1GVywu+kDbBwmYdWYlhtTlMmuTpukws+Oh7rMnIpiKLqNNicmG8hZpXwpDSUmMDiGMrbW
4Vo4WYIBCHfN1Ji2QsL+6JSRS6ajkAtsHyWLdMzF/gqOkb9/vQfpICctu8Y1D5IUXHpkWYs51rNY
GGjNsAmO5FzwhTsSvg4Fl6dz9w6CP2kLYyK8sXyPrHsiW4Iv2vbBGCkY7HRWYCPiXSMRRx6MF8fr
T6OZAi+nI2cOrA1Xx6GZrHi8BluP0yBLhiXc1iF54jpU/fp2isGFO7m/fh3OYWpOUwl9mZ9gc96L
TV0bRLFqp4liBBHImSmTgGlCVrRr/pPc3uGbh4Kbv2T93VI4oWd9ML1ZYz4zFkE4atu/12TdKLlj
q3VSnoz06906QJCDG7mPgJ6hF56yD9Bc6uMaFnMCKBkkHMNgZz+aDae+OWMr7appU19qb/n0GuRE
1ETLN7wHl5ugTOQI4khQC7hKylFMTKge/HgNrD7MmV9jo6SxDoG+//DUxln9xswdv3hI9pDno6AF
SV1xBBP2J3UehjAVNkipAIsNdNsCkd1wDFrJiwaBADVQdu6wIruK4Z9O7q65H8GG34LHGlXE+waH
t91HGprHKloTFHeLeXmRgv31cSN1dfxb9ZipWm8xX/+oaczfsXkX225NCtV2pg7R+CmcTPhE5IQR
cgNjtiVoiOYIP0JYIQQJiMMR6QFQvSnjO6gde5zVeCklTNPi2GzNKSjOGe0HfF3hOTMPfnANS9++
Ry1wy8o5GNeWWswSfXNFrdA1zmCo13JSgh2VTKI2XxloaUg5I7ZruDKleYb5SRPCLeaEwkASKPsS
pzezft6v3g1MQ86Tzm2B0xdHnNhxMTeU4VLRwpklFVp8gtZJgTZrCSAD3czDMFNlUbZwRCxc2gtZ
BAxTmNSEPU5JsP+bu5wr4vmUa2v5mmIJVe83ZT8/SRljxoYkN9RlKOgKs5MZ9CuV7GyxMrYaekdi
WVP5RkHmkoVLKgFaKDWYai9GuT+JfE2reCGe5WcfprbqILPGmWVQplFXkmyRZ4SIo3+Q5GEPZk+2
Z/2k/A5LvSgqs4ShVgwK81pZww98DiuQ/pBqXQ0M6zIo++uHMGRSnC+fbKadUx2BZvwPPViuPaCY
8uyPjoeX225FJCVEiEz/zMUGQrf1TJZoqznF+arMrtAHQIGp7VPNuaes0cWDITAWTxZhkzPbDtwF
i3IrbgC+Pi+ZuB3LtfgZB3CYfJF0OVCoO+es3H7jkOfApEqlyBj/IxRlJ8M1/YXhYfRD9JZ6CE+1
dlwZppT48DuZXvLrTF4tyKg9ZoVUWTuN8XyKazK7Vp+XkQt5SpiGvbwWx4wbsY/r30uyUkQPGWIk
KGNVYDGHE+B2xCsPs3W9nkZfLh7choThB1dKPMnNKb8qitjXHiJGl9RZvIWMdtcynImXRtjmn2IL
5rHOz7kVC9gaSEBnUxFHMCAKcr8bpSOkTbmKXIn9WBu4fJh11I9xQFdFYFhYnvxbC/TR8PCWB8Bz
nGDT6E85ysCCHnYIGQSHOm6PHqDmIVt5kwu32AoVYWU6RtmVBMICr/dln5by6H7D6XnZ69LdfywG
445dWgKIlxKTwL6yP/y+mbzREd9fQsqxFluZFw+oqeZ2UTdqZ7boLybEm4NZ0rcAO+O1A78ZzPBi
rOGmTdFRmL6NymwEE7idWTOnu6bzho8nMVoYM5Wnz0Sn8q0K6jrsHeK2k46IrgXN1U+NmvYCa4h6
8/9SF0ciik1pkwtpbzpXq1iI4RPSrRqL1ozWBgpvCYyluf+qRA5T4foPbuesZIvXGS+Y5bclrDYq
tBmpKV/a7YyKrNbOrdBoiGTuOXRWduFUNO8Oe5P5T6DbQ+boSOmRF2GfleUkiedqQIjpZN4XzS4C
aQQonyFi3/xDq/Fg9lednP6u1X8fowoTqocMs6e3CFnNYvOc8sWfcTQMIs3Q7I9KhwF9cid2A4rq
UtZxqjwmQsjFNwRxm8UcPQibpeGBKO5UjqPp/p/Lw9lHCXSjP78OnkNNs9OjQ54YA2j09TkDx657
2+IbwECL5c2Us2V13NxoiMAma3eFIt1k9oBgt+G4yMg/gyNWoT3AJK2Bqqxe5uYD5sBCBaniF/fk
O9qogGQewIdoP8Z9u9GRbgGybE3tpEmXHPwTagWHQDXedgRwlsWLJIr/YwTlL4xiJsox10GizEno
PNP+SwSEpHPZgH8MDTKh7yqXDsgIfyD24DlOAfXX05bV0ORnjZMr37822RaJoJm2F+Qcn6G0Q9Vz
2xg+IefV0R5sLh251A/JTolMKyxzbnJdrM80yYFJT+zXJfxhdZ3fH4hGRfjgHTd14rdqWUTOjiU2
7qd30MyKGaRtUDEqNvDde//y7QUwHDkrQqCI7e15uoWnoGvWYEeScH7GtPD4pFPll769v5iURzeH
i1hyDYUKbaLBrXSPUg3d3oykd+XKPZJQCAtacTPuPo9ZLa19yT7V5BI6TDNV/Foir3yyz13n6CbC
ROxqKb+NzGiUSSkNl4UhYBxJFpEs1zshKjA8yo6EyMgT0vM6TXHaR4Su69EpebCaoJy0YuUEagmp
S0ePfxPucB+8l2pbrM9ofVjribYlai5R12N9B0ZAU/U0L18H8rs7JKDTZKknsp7eR0arK89LU2me
MYVgwec8Sd/2DNWjkhwS8gFHnPEZEq0qDPMvfJV877AEjXowntx/R3c6rh3233kqaE0VCUi7bPOH
s2TZI20bvjEUqU/JbXcaG7OZEyr857+PgNKaFZ064aDbcWWHrGiYg/JmW45U/AAwoQFNy4qnQ+I5
1RAaakplHuXsPc6kpTda0imKIOZHAWvfUSE3esqUH23vX41KfOfC9kTNvMpBGsBrwfEepfw1GUMJ
32Jf4B7eCrcZwgJP/K1AXUWlgY+2F0mbe5wlDRRK+fq1vQdGpKJ1m+Mcz+l0ZjZ8LSfOU5Xxf7R1
QJHtrZ4AvxkhL+7l5/ceTJ0UKZ/39jZJFXw9JpCm1Fw0lBbeKLA+zN6h3xDZ9eQgxDLcxWgXOE7+
1iCJBbgML8iBiZL8FJAgd+3lpcfqI2sVwT9PghVljIBg9g9/HlyKheOxphXBpiNfxY1OkH8hwC1y
8Eggkel6Q/OE6ndCISrLXOyqoxfHA0pR0QsdyizRCa6aMXFEs6vgTPMbAisF8S+4WATyiyI1jYrs
yWCJ5kS1cjPFJrKAxpAKy3it51YG/p/j4QETa7dIJb0KlTHU2+VHSw/e3mUXqEnxXJo6lcpyPb3w
ksQ420CO/oWkxUihUkgU4CLx08vHR0oRBizV5VuXf7gXl18FnpIW74XPqlikIA385ZHkRtv2xk9F
ZFgOQK1ixhM7ypaO/sCrrfjA/ZLY3k1MNNtQvSdJFScIHkZefg5HEI1wej0u0d880LnztjszlFOP
GuSRRDYzClQsNsiP7jxcH/3VzDVenNLiS0Ox3LJx7sJifzcFuGJL2fGYxLMhiklThy3bjSuhALtH
1ZDuzUz8prhDf9Qp5DFdrhwvaFnWdHOyKMmU80Vih4UdLN4mx7OuLMQnshNyB62hLyndhBUH49Mw
vgX9nOzT8dIc6mLZj8DhoaNBWO8q8TFl1IUrrbtKfOy8ao5eur9yAissN9EUX317IN/TMJdWp/GQ
R2uwYYpCsuMp8OySI28iK4O9paPnDMjimLWJkzBE7DJr4CQjogV+Q0kdaVc7ToqRZ2juLAeGXKhA
aI3M+bFWRtgysUtS8+YwbiTOjhTDvCFLlFBi2gLgH011PY7ONgseni8baxuqvZg7rlnj3iruj4nt
kOpDbvLy04nwJ8QPIRAXk+f4OyxHW+7fCWO0VqO6fDjECS15HJnl8K7h5S19JVg0tWsN7ZFJDhM9
gKkgEHMpXdBxpeExbqOG3iFmgt2xk/XIZl58aOUXCQPcDZswu1TBCReYRFbqOJ/IWnq6Zgp+Q3RH
h/uUlBOsgRWlgmpsGL/Ahdug/ia4EUvSKq9YIBWIUmk35ERp0h0FNdx72Hw6APRJ4sAZIxEECU4r
doxEMoWqa6xEJyYAH/OOpYtM3HrWjb+lRpMUdP0/hHRUenXfe19BWyG5v57sfVh1XNLsm0oAok9c
shXMTzbqTZ/nbcxLbb6hk11aenjY66Hkpgcnp1fNp31qu4GswSkHT7LsK7+b7iDNEpgm8Xn302Wr
KHziCLT6Zs2P1Hk2HtOj3DJMM6xJ6SgCrmqicZigF6tMlbaa/bSyorPCFz83PHGG968ptM1yLRnI
/4966w01H5nuTZGRiPoT686Lid7jJno9hFJnolol8tOUlxTFPHTssqOtf4qhDQSKkTQjPv2yNtRK
Vz0hX3IrDUtQ31TdpEodj2wgJGiOj0QnJAxyu4r1RuXhQeit0wGLaWaCazIZDZsTLJw03meJ/EQ2
Dj8NBhmrd1gqo8mhfM/MmUuLTReFVWn7bHeuOaFW4y+R6iLqXWJocrNC4dXvbbs8mr/U7PWGN8Ne
PdfFxRzznWJgwPw9qjMG/1rbkvHDbZxaYrOOJf9Tdfmin1kxFFsk8r0auHPznEYH1xMTTp9LkPrc
Vx0LKtjmXX7/Swg+TQMPibPPH2tPIGicdgx+h2FS9ZcOUxHSvZ3GSlykHAq/b52MrSoWnUkcAY3v
SK08ljE1lVk+uPJK6fycEVDkvWZhIfOmfcGML8bUp0cspaJ4VFU3HKG6bY5Lb/Mv2ua1FQlRjHk1
VJ0rrDYjJ0GIUNGZ1wujYrtNmusvkxZtAv0IUej/JoqsceXS8M1s7joKtTTlBy1i5T23/IboMgsX
0we8xZ1RTjVC2NHKfVY0JmkO4UNDXQJCwPRPUNdDmaRUV4ppor2hrTus7CXckH4R8NwwlBoBwuhG
iCaiIiveYDoA1WHhZSEanBF9c7mTRcJ4Kf9QbauU1j8Ft6qgRde/tbmtdNsFdfpxGMWLDbyHT6dX
LYGXoUeQX7gA4WHUzUPuKb7NWclfHSw7Gc/9w1R1V64cl6xF/bEJpghRUJLXYORNwjULXeh/YTa6
0bHGoIH1GDYvUFyQT1kY9jyBjKF05Uca4yAsCT2h5J1biHjtxulTednIM5wnFTPOGe/fdF3Ay9ED
jMf07fZrvSbCb+7WG4Nxavr9fbOL7g+c7JOqheYcKgZoIGPlhzNHmn7F+Scq0oUmZcntgOl4Gbrm
lA6Fl3b1Qu9FOYOBEXAW11lFIs+Wplf5uXaOnWH4EHIulNSQ4kzVDcocI0NzcPzj6rE821I8dV7e
zPtesRD6aE6La07NENpWleguDUTzYQLefW4u0Jn2nWmtNs98YmFU5MNN9pIwlqB9GoYWiKswG4fP
42n5O7ZxYXAY1qime8rOba4PS0vFYz1zy9fcEAoy8YV2VgroaZapj2vSaxNcTlLj3OfPfGy6Hu3B
SiSzY4fBUKI3N73XjjodE5P90KBLK+WQK90Shdeo66qdRD5FS4VuaQvCkY35zQM2+45FmttzD67r
zuV4u+EmJjYR84c77wa81MWy8K+hn/lGPfH9TdEx7BnrjH+Up63phV9s9AaIfINRWhO9fygClKSB
A88d5aLGB0uspqY8pVXuHR8I3XNaE2uo7fzfpaLirCFykD3hBHNZrhAa7QQzqyiHTnEn2Yz4rVRJ
Zowrn1r6HUSlRo3BmO9o0qx7nBzTbsjjkE/fxmf0feXN9MUKrfIHypcQG4adbeJGSkmGxNoEzxJf
4QObI8VCf+fms9o5oZXIdmZxLNo3JTzcJdnsQY4U650mfADEW2qkbcAHKy1360U5rNxVj6ZN5En6
cGtHgaLPepSFp0LxTgA4FFCHGNOnFiuMPk6Wv2kYZ5W83o78R5Dyr96mbXLEUEsA3pwmDZ+cLDZf
drv+0BHlUdKnNmTZ3rTVdx9O3lRlc4wyqSGQ7zo+TnHcDpoVyafTi237w8J0Ik2A+rfQB+61N1Ya
EhvOMLeOxCDpy/dGKj/M91+A/ykkBRO7LYu/KhMB1IUsyDMv9nYU9DW1QktWIc4/X8YeI07pN3k1
mJdBFSW65CzGRnUk0pgsYaxz7TX4F6DH5CTmq44ESDQuMZS5pdkxrwopme3ykNH0MLbgf7exHU5k
4IXMIzlgTAGjILKBdSADgDZUbXUeHgwyRx1xhwvQBvM7dSFQDYJfNLeBNvv2L1qFKpadfT2bgxgY
mrL0AUkd1i0lrqjpE4n/5Iz6IlA9/kxMbP/7Cdt/lVEfWvhxwYkPy9XxiA0WReu/z4EQcJVvT8t4
xMQ+3WEoYetMUUAvEkuMUyLXp83bl1YG6CmX+Aa04EiVKx9L0fNN1R1/6RHrwnnavkMa3TjM+tJO
cykHwePJ9IBec0EcrE3kYjdDztJqjncP9e3mssVWemo5jDa60nyHESetETjmAVhCC8qyOAX6Xio9
20oU0iewJIlKAd4sDz9CG6yLFJKtEZ5Uv3B9CBj9qp3YPj/e/cDLS7DLyb9xUSRts1NepSekZ+lO
N3gNWM8QBkgpmlLCXhyn7o8a/tE5NBNR8qH/A4B5GuS85TWIlBgtB5Yg4YfAbWmcnS9b6rNuTJgC
qXB1bS4sqYOqpItTr60UPc6U3E9PJ1rUdMuIf7ka5728VmEscfnElKVO0LFSf7fpJwHsnfBOqH2w
SszL/Vhr7eNs/colznDYvUJN6Tcin0CgkHgyuk1ySRlPmgovmkimDTpTc0ib/vgA6NH7tGr//Grx
9ZjwY52wB3pWpmUCrwfMceHzxhlg3PZOwYyJ2l2+Fmlx/zqoJxerkErFqIkaIN7rmC59cVXweiVa
xo1N6WQfqpBO2i7gwa1E2+05ZuOvthz7MaiK0Fqqrt5rys0xwW0Aw1UFmLhtUcy76S0CizOKHE/v
qDQAA9bpOjHelm53m4AcvYqk2nChxWqO1jLgQzQQl9280jyJcfUtSgrwxwtz8KpiSC3myp2YuUKw
s6fK9w68gsNnDPO74YuXpUfiA51t/kSvM1pTjdjtY3WzX9yzZWE5E9p46CMbia0in/GAnZhpZGiG
C5U33kbeUdlh8Lmr4jDnJoj76w4TYjzAqqSQCBP1psm1Egg+s982rzlpPitD1xpY2SDjNqhmVzaP
6e70IILVzaJV2D83Qlk9hIB6jDlkGiuNoAd9/34UwIb2jrEZ4FSv+64BQiJV3O3X6S7uASkhWHLj
A1s990UqMbfWImCFwlc7ZzgFcPp5ek22re6xJd7Z5m+44p6KItoKiNumqQ802fhzL6H7b+l1shdW
ul0nRqmIouf6AnRFy1mDRJFMz8s/6D6XDzi3XATSG/b6vP2IeV9yE/OT77z0Vzw/dW2yKvRt7TbY
K3luiy2KjtXVeoqXgTchQzIBqp7X82dw4MbXWvVSHaYnRZIDSaT1n6k2BO0MJgB5m9HPmBapmj9R
qA2oSe8N5bguZd8gx9TGGMzPBKGlsEi4bDY4FyFBonqBW8e6+ARoMWqm+UXA0zoEvqKEEtHwQ+kf
aGSYVsO+M/SqZQ46X5CCnGidY8NkE3+tnJVzEa+C8/U0orKbepIYeV9VSpbOPUAPcMojZapvI5cj
jzzv3nlClEMeNBEKql75cMfbJa3qetlPdqE+p9p0S7USbduRbuAN9YXbP0axl3bQV+iWb2d9mi4G
helUliEg4wHw6gmZQL51O3CWzW72lIBpcYEcKv7dOgKlQJiWV1Wk+neXElTVqLuUa7hOQjSWjdR+
Q+20ttYFUiAP9HMCJgsqqEhNLRatTLVobvX4GHvdVsZCzIz0JtA7wQetFXxdVTiU9AXcn1B/sSOk
fMT+v16sRusBK+wTReXAnfb4LCoJaXRf2cKKgRAnpVRK+90PBfCTHJY6oKUiFGpXsV0OLg2wo0wN
gfZLSkkav3n/68FJ5LV0BBzSK1HCEz+dZvEfqQOWg+0DNUAGntg42w1HbfIJgO0IdujZuhEHquZS
xoWSS2WoIGc6nHh6btGdJfis82nTmAv5X3BHqp5/b+UNVO42Clk4tkjxl9tE50Ab9R8ypg+mAp7G
1qe0SkNjHlhGHPjnfKpx3+aGvFqWUgKARJu1kywFKnhayrKfjA6FqdEr4AHSfxAAmBVHKAFz8L3d
loyddcAcvPTnaS9Gu6/i/icTsMdSEMvCljbzZgeNFROhKIqfvuWIxKiVSFYTcHIZqTiqMXM0mwnh
ZoXM95ET8GO1npXls4ygB7xsB4ch+T6t7y1oZQj4RU8ygmI1Mg4TU01YF8lflThDOwQc+GBsFLC7
xUed/6yU7WVJsPrCvjI3njrFcvrUc02NfRlbdxiOTm0hn0ZNnw8KZTK+SpcTbmTBKUhKqO6xYEbc
HYWMB+zQZ/enCXsbZMJ6fNehziy0N/YfjLqDg7wFXqaCeiR+tms3nuYXbtyzVUUJLqGWl1RYUgsv
Jneu+wxXvpITOoIRx8V1Tf0tXFB2QS34X/PsectYeDqCMRgWsR+apHClRi06FWHCfuvwyNL4ASg6
m6RXXADMazxpqhuROmEMrvIxMQIn6PmJRjZDS0wsPEGXqk5JMIqSDlo6RJ5EGL37PIlUaDwnKYxZ
/ZR0nH6/En99YQDLxNXVeO14Bklc9tcffoovBOX16e1nnWyRDzzVlhisWAySHidYBkrPffzyXx3U
gvppsiXtCSAJkNf7J1OjLp2PfyExBoQNtoKQp5eGH+/5ljrs4qTsjImWy/JkRGxyOC2fhFm1azwT
sR14EDaqdDOTC1QwMh2VqRJ7yaVVMOmRcWRv/z/8m69uteAUnA3T68C7t9Hi6iyb46FJiMTgwiQj
0XqIRCu90F0mtCxgSCwBH3T4AYrAbWLocjxOBDZGBD1vaUlG9H/UkyQRN2txruh19xXt/AfCFyKW
c8FD/tf9d9xzGr9JfdAzGZ53+fgtku8nJPk54jDEBZeGyKpjgIR5kA0RfkpwAHl1jENqa0QjCugp
F63u5A8XRKkJgiQ38OLz8c+2m3U6J1uGcgx8ge8vsc9tVpbLAbBmb4qqpds0ik+SU99o2mCQjDx7
WlQIH1179BMt0kBjsS5IITxIo9GavpqXW9aEy/mU8acGt7LvALK17xHc3RuWG1koT3BjWBAQA9OZ
7jwwWzRMVqAtrcH+ZQ/CUykfVn9v4eqcAVd/N0+O+Ntm1s8FIIHqfBJqA507WYFcffs4fXoDkj0H
RK8laOYhptdOPef6RwVYHX6zcdIO+v/zHHrxWet6Hv7JBJpCMfFl/tp+fYsJxk05+DNNZYHheXjz
c51csTShv6tbCVTsO8M8fg3i67a/jAfg7fRZNWryDHVruaK6t17LR7W7kd+rndmwOKbvRrxThmRC
q8ZWijltePNox5pKdlGkRWgKtS/5LkQfQw8QILTx1nK7zTDqJSUDEV/kzt8ciQ5njI4OKQKbjwl6
1rZLDs3mnBBQNLZzCC9Yserxxqbdsrc5DAnuTqkqozibO7pKeLQh95kaf6gkzow9ONLsF6sAtEOi
rUz0IoD99Uyvd5ehFntg/12jDRDPG3ystAJeBkYYDiJXh92sF72iIBf9IuZ91NtseHG26o7uFJoP
BenD1T2bimwXauTx/nbbwVMd25XDbLpfSJs/2Jb0j5MTJIAHwkY7Kc0C0BSicJHCboOsIBXPKnWM
mcksubAmkiOk0ckWXMZtSrje4W+8pB3s+FD2Sc3tpPR6qm8CRStf90X04kbgbGh+sKHt2LTBOCIR
SQ1CdvwHHgIf0zdOT3okzhftqKHP0YyDe9znjzqTzkOwXUh8DZjEe6HnRVuRlT8ruQeulbOktojQ
yT1JVDF8fTkiWGtYPVIEwVlKgtmuawGfo+bCFsrUEVGwJAJajd5D9nSdjq9yzLf0WnzPRMLdE/Sc
iPuB0uoPCbj+q1SUIvuyfPT7QDZNQbIquLemEcPTyVDF4qOBJO3ssZG/A2FKmEtc0z7c6p/FyY7T
HoX9e3tpcSJfz4j0oylNR/1ST/uzA8VxgAL7ntFJURWDiDBvQj7l96+M7HFMSlL5teaRlNmuLp3y
HbDH58uYy5G47CNUwNIIRC/+ZetFxY5WH9f7Y8Nl3G31aD6M4xU1bej0MAVqb05ZOCZzsxcjHUWg
gRTnJ9Hi/CVttPkD6gtT5kmxSGhIXGpykZaNSAJO2GbQGuxIBxYS9JQcHsDTbCQ/UMCR9CesyTAh
Y0mqAeAq6xn/EOb332OD7DRaA+6Q+UYrGBKK5/o6goi3f3/2d/T4RMgIR6Xim2Fs7E/ErADUEQ/t
anh4Nd3AbJWi/La1HUrzurQgis9ck5DAf+yT7g4XOiGWafEE49O/xGeTPXIvY84joIA++ucDED9r
8s/7VluPIdBozfq8abekRbAU7th+e+NAP+LbKCPBIzqZuyKpcvj3k1CiUPxi3lEFjhlDnoMWYLqV
UF7PF8M+1ZrbtcPGS9haws8RJc6S88iJRHKheXaFCLAE017uPTIx6W0r2B1d65pT9J875oO+a5Ah
BYZfvbn6TC6hEmW6hmsprEllqmF/bwNoGOv1zmMWPxqNNm/nCZq7j+YO++X8qJ9tSLWngTxcL80k
ylJxRc8WWc9wh7JmE31hlb6GzEwJXN2fmFYzVnNYnvE/An5U5FRa5cWXQ9deLOFrbCH+NLBP6KRA
x/9jQL/vhQckpSWP/GeNXF/dvN1kNkE7XYNtqTgYjC3KV+3P8HCjORCUAHWeO3CCz1EFPkZCtJUE
OKmO2non3+blL1mvgbfG6Ei+b9zjbM3KJaptwY7ORIfhAIjBlvnAg20XHndVp2AJOxMKjHyBm5RE
TqD2p9wS/cwwMoZ9uq2Fgmq1Zl2mHcv+VcEmwXIavmo8QfZy2vMEAGh0W/hCF4pLsDoddls/dxNK
lumx0MOHcU87PBujWlGckst1HStFeHJrNCJN+2grbMyxeY0kxPx3zrUN84asRqc1mpPzRFaVdOL4
NkFBeftiuPWmlk/7IV253dzFUg4tjBtILHUWNRX+3vwkLYH2/P54L/Nrsj3Qz8jP60nJozZdpe2e
46aeMd9FfSb4JOeXytA9sEaZT7JX9eU1ej/x36QqOE+FML9wFyhOLNzoAzxcAiqyt0VgHdO7PITR
GdQ9e/cGdUS4JDr11hLlpBCzqDCqlXH9539DyiQ2T8wzCD6cdaryh7yWCLbuEpyWVC3j5Tp8IRzw
JxBpF6saeYKGSRXS+hwf+DZVobXd1GFk9IcI+sEeUbKRn3Xil5DAvtMF269KY2Who27DuXqSOvMe
2rMJSrKrPgHBTN9jXC9XVShIksUnRUdKILZe+GRgdHfjV2OLd0sOVOjqJTmDXNuy3CLPfyzIut/C
r5MPrD9DeQsBP6c76szuTE1TEsQB0tSwkMtLzKtxTm5leFfJ30PdoI1v8ayZAd0scjdvT/8HenkP
GyIpjyaXEuD/CNmHmhZGlPg1xFbNgPZFNm2ddWGDyOczSRfyQ6NIAIKcihDxO9NTqC8WkJT6UxRr
APO0pMqbD6UsWIDg00xukeiGvptphjFk3Mc/PD36eUhfr+ldANfnBUKmdlyOguj1gwUmSZU7VZef
emW5kKHBvbbwwoHZz/ETt9COV5U9pNgzAuFC3LX6RaAbm4boPcFkRGawog20Hs7C/+v9rhRnb8Dm
LlIeWY73cT7Y83/2bFhYjO/BbEY2etA9J1OvN+DtDPosueTwBFjMFWmttVfpZeWb+TfnWyg0QZCO
lcYIgZYn8RbkSyCiigtGJNRkWMKdSoXAd+Ranlxn7MgJ5Y/eA35M15BXMWsHZmy3tQTLWKghZNfh
ILkQ+v2xdUkEJBqkYXP3AqWfCmBmXHavX7Vg7XQP6vnb+bl0Wt5lo725rl9dDXbHjr9EARE0Etcs
imoELrADLdgiu85zc0e4tXOkP2myS/SszcckimXvqj/RRtfSAFMOYTTPL+/hT7q+n0u+Ja5KxI66
1RA7OIECnVbnO6QjR6wWuJg4SlAHoJmBVlptuMY1nHMwp3RlipWBPimI8UGYpinmlf/ydyMrWvgg
kN8FxbfBIq5YEV+vehTUFX7j26bA7RghQz24Rvj1Yka+KQQRfGuzZdzOuk2m1mjyPQimkgPtKEtx
veDJTG2X5mK5sPGjC3JSL4Db6B8OoYflCIaFsnJgstm6YYVoLw9VLmry6p6bjFkMQjT64IF55cn7
Rq3340Z3iS8MPzt3Lm6p8jhqsiXjnYj7HemLdV7+hXWEpuuUpy8QYXhU+yfrpRk0jjvM9ZBgIqXJ
Zu5XgUcRElcoNnXXIw8WdT7fnfhanbB8H8WUlmqX3SjqXza+OO1q5/ZwK14G3hsjhJd7aHNjq2gm
wDOuQFpDw1RWznkNWUa1K4o3f3gm91DPe8gcbhC2w1wU8PZnu44wFILd3cemXI6NAuDJICkM6vpr
BtK7exvlQP5iCR5UKUQp7F6xl6sofoFQrmabc6CuoobMA4/wJa1jdTzWMFNEqlWASo5QVThO9B0v
rM0UYN2VNNGAjXp3YqBMLYRMWJEnUUnHyb82CVbgfOQ8PoVDuUE8HdiRpGb2KI9rMvDhn4foW/Ly
u+vG0dtdTRnt7e0xXd/5lpknAOGPQhbBqUXW/mdZmHs16tPJ9wY5QJ6VakQu7THOdObw14+Qu4sz
m1ou8zLEV2wO9ElrfUtz4BImohTh/gnvP/UxT2a32sfp/reua9kI0FPVgyk6Z6/hLYfDvayOiVdd
jnOoUaxIrQSBFJGXL6DZgvLZsuDd9CdX+LcCIWRz/toHwuBcgVWZD1SZHNrKAPMeyY5Ih/H4I3V0
JOliiNZLd65/gi/OUvawN30u5wr15qRWsHBYVnqd2oNL2R9aNdH+dg62Udc2+xm/luJI6qn0L2i4
5kcoUc9eZZ94mfX7n0oQ8QmpKywQWBXPASG7AZBhI/h+8Jfw0yvTaOV5pSSLQjTKx7/dB+TZcVto
S23UHGEEhTGgPCRmsXQ795Em2GOT/gn0dUSZkEMvjZAT7t/wS/8jWBDDUx+i6TJ72SWaKX7FRCZa
RvQvkIX/w+1QJ8D96xgqQyqA6fy59pH3OzaTlbbkPZkk+sRzmy0XQRzEIc+mxWdA+dp48GvGvoi6
aNzSbwCs2lZShuzQ9mlEfCPWxdM45DWWcJdpdoQSmME84AKhbV/HnP1G5oSZ/vsNP9WEogS2X/Hb
KJnOQqZhybGXyLFbChUMDrB0JtCGK5Dh5fBY4HvjDN52B8VmRgPnt1Vg/tIKDJHESsGVZV/qnSrt
KwYjJDFR5pSoAMB9cBYQJYLa54Po1/Il7IW4QzoQgnNGNOSQRkqwuiHewxnfmAFrPVMqSzpZ/BqN
OjTNzwCRYTdiYRglO9RFJmrr2XNGVSRc4fKt3+MSkpT7QikalwVtTR1e/UQ1//Ljdcbx0dlsP5U5
yqt8BYoPWtmGsp2huRtjLA6MTdrDVnkKHKbzFDuuhTcB2v+iK+uXhe2i+Uf6TXTzh1D/2yOJ/LAZ
ejPRMjJ/HFlTyPuLRjoUp8Q3PjxumH6AGL7fByHoNP9P0v31ffXsdedVE4bstSyBT9Ckyouw81a1
Swf0+VQVAr3UpfPg0O/OqPy98ILPfXMDjNddgx+4yoamkZshp9rgHaWh5wfkHH4lZOHt68wRIUzB
RgRK6mfoV3SVE1i4rnALl2rTidoOPm6101oEpAZWhMAshA6H+aYmBhqPbwYHYirMwSsFeXXgerF8
JUga7djEUIyY3aVQaJVRyZxK+XWi2HUMpaNRL7mljx2OaWZOMOvqwXYTLVl70CD37v8qxqDBnu+W
E8qJoPaGSbR1cOVDmtb9Pz8X76g8VRPpeYdHHJKu5xgOFT7dCP8VcZIes+l7kYlN8wikcpcu/emA
Jh2XHvjNT1f0qJGKJObtpqURUGh9LMyi5NQzC1l2R/SPM7NSVXtPKjnvsXz0AmqEIJFHw2+8tL7l
wCXocqlsY/lISfNxbxAurdzYj1y0GvP5Rh3oQUhP/4whnLEindAkTXQLA4AJ33090RKpse+xGkZ2
MNnRMIof1taDaAyPnDpjJ2AbxcXFmRwKPQMjQs4dfJTXPNIb2XZJjHIK+3ONCXAivbhRAqLzAVLD
5fc9rkQfIbM+LxGZrXKay6Ye62IX15eW5JRIfpn/lpoQVO2HhSikBhv7c5/DBnqojeBa7tY0Pfat
ART5LR+PZ5jSmAw9u07PslIBtt19ufTE1pxo5Ptdj6JmQtPArUYHCJZafRUPydjLVtlXpQgaaUr/
pFrSy0Dbqe2NvEYavGUoM2WPfUKJWjJB2xjcq8cfYedK0+U5nuJUjoQiKZjRWilrrsZpO1rTHwCH
7fbATZjUN9oAbPcEK2IR94YQF3obrA0s41Q8Pj8dNhwyzww2Wp52QwernmJGPI/agfFJjOApgO1K
73V6OmpdlyZqFlQVW4AvO+ECU/3YMnOzw5kPqa+r3G9BivzEz4FtQ3N31ohszNzYJxlI8BB+IJ7Z
LvMQQcjN9KECpL+3pFzLC75KSSvrAhizgwGTjl8jU7okOpACpV1LdbJO86upprus6UgkG1n9qtfP
BVVkhWeQaKfOqj1l6jLW0Z7HWTg9YYNfg96TD3uGgYDV+ZJTyFpHxAdZHm7ew1rkgnAfPJ+Ukfdi
0tndjJXSjAAwmlIclY3yULw3F6coIZQvCv7R/GzNo/bTsUZ7J8m2WQ7JXCroBh6MnvBtXJ10fqxE
PrqtMQhs2bm8UHh0isLc9OCLTLOfC8autTjHDo7ighfHm9K6siflxPFsFQmdzajLWvf7msIVhI1u
9mBOPN/rTMdfCDr+OYjY+ZBrwSFCMhFWxGGDFY+0IG/eEs63eQx5rQSpp9qu7RCzriw0Zmlyv156
qPZQnEjMcmJGZ1qlHu7k4Ma7FNQJo6VzNgtO8LKTNQQB8l/+arEyE7Ird8PSVQpI/6aFq8qurIkp
advCFP6LbW0X3k5N0655z4iTKjrwLI3uvHfDb3z/fP5lGhhS2N2bmDPrOb5V4j2h7Bppqloc/WoZ
5z1BHU+w+7fv1lOmdw1EVbRWcG75yXF7HkGURRPxZF7jKr0W91Dq6YuUI+Wz4iIyRybW6RH534tD
LC0D0UJUjiyK3zlYCSEmdAsis9bQ83BqLJCBMiZTNexh52FJ/TVUX9w8MC57eD/Lh6iaN/lQyklv
uu9XPA+dXzo0/CdVpaO2diLNlh7nvuPmbrcnn09hFuNgfizNK6IBns7vjSoRSrCksDMw0ZF4dqIl
tMcTLkPQYFTRLt5/+3+bqFOmRppr4WM95pSW2GpJeRbaxYdWTsAYgx5xvQMv6NVJFi1pWtCLcKO0
jDux1f7mWT/eRCOKSJF5hMdUuFDMEkuVk2xDkBd+NEWfTTjNVXXG383p6RafNTv7/e76OFlP36xV
oGnvwc93eXjBf6dvnC75t5Vpe2VL73SLO46+GgEefPYloiIzlTmv21lCvahvJjyXK/13fO9pYyy5
+r7gkQk5GviHziRHtb8nyvSaAaKbpJKHz6RRZbN/eC4kAhY58DtBKtiLlD6T/M3scGEYQZEUHEQf
VhFG8ApcwcpA+MPpjg1zxZV3KXx2oznDZuR/7p0R8UE/TxluuE1b8bf4uR/wJnx+S8aCZ4gtUgR4
Z/kCRPXvW+viF65+kgcV7yiXz5s9J2bKFdMPUoLU931gl6WpY1DZ8QuAFeTZBRQfOL2D2hVJjeIy
pkGl0OamZV2AoAk0qBWVg0P/eJFQ7kdQHbcYlO809FYwbjRY+WBbmEkHJCOcz9EFSEelPeZjsThd
+mcsrdFdy4PgtQ2/lyTtpM4Zyw5hx7kIn5lhSLJNRfVGyGmsChWOjg09/rNzOMRwTVXfoP+c3BZA
GlfjY0ENNrmS/4EciuisA/tiGdXiqF1D1eT9L7XrKOaEPYb+pC8UEDoq7IJfhdlPDfLwFOMIfMvE
r6gKsQfU/bCvD0aS4DZfpL57HxDB/oS4Lsy9igxkSirFmRTVtwZ6dEgqKY99CREs/+ZfIMasARoP
fqKN0C4znogS+W1cyaCcdSs9kF1dFSkgelVKs03CLq/GHzgu/9Ld6323qfna6z97m7UgqmPtLqvl
vVaseacQ6XB4rKHorxwPPnPF31aMMvhPOE8oaHPwNk0kx5Bqk3Qv30k6tPp+KkUknVTbZDWDLKTT
TL1HqEFMiU8fg7lswVkULBJ5st7RU40nVT644Cu4l9bRPZe4dUXbDinZFGJ7eDZcjqbC+IhYpRF7
zPgIs6XGo5Ko24mMyaAVJISicFhbFqcQAnoN1lmYN56OWwJZGpn4srHXeF2sVHjycSHLYK0i3HW2
ZvlQHS4iknUKgnkh2gEqg8W3XExrrmgXFM1V8DTgf2FYl2aMlq5zk9Vurjz9GlRM5sVuxM60rvfy
fymHyfulF5g1qu1A2VEE7VyeDT3QrJougskScsxsjdVYEVxvpIBsxBY9HMbqX4JnMdDXmR4pc2rL
TSKm6MA9moHaNRD+7VoQP2fPqo/3jQ966XTUUQUz2+YDaongQD6Sa2NPEXIGSiPp/Xri636g4/cx
jthW6Vc/iQ9+7eU4BR4jM2gVFC9owrrZ561uovG7ereGveJzaCx+jC3Xqej84A0juxS4tbWzcya5
loMdsviNzCh/D3AXue8L70Rqi4Z0PCatZc4CNFlGsDN8WSiBrZqQ9M5ki/9R4Q4LVNLvvAayJ+sM
lXGkRQF3mdIJWS5oqp3NccO5eurHYUYNevF6RdbZ4cDbNpMb42ydW8U+8WLVeVVZwa4E4KWvRBKR
XszAdhpwTNYddpo4JX2vO2/npCsgghq8YM/Ta1YK5mB771oyCbHjNEJ76d1J2Sf2G6PycZKVl7kk
3u3eCejl4rh3SINt1VWpsH7eZn/Fzr/HHYnMd+TTkD63ASNA9KQgoRWdRistOlLTkisIJ+i9WeGu
Vj+mYxPCLaKdv2vzMemu3XJN8Nhuu0hVIAscv5k2JCS6yP3oFNdc2LnltYc2Pu11wslp9fcGJAwf
tR2OoGN4W5x2o1QzTIXyRumT/o/R8O0pMWUiWjQ/V2dpLsf7smqFbeSmf45cdKl72Yjg1B66H97M
ZL4viPdXeN2lq8y/GqjwvN6BWbskDBpqOxWOddMnCPWWx4Uva1QdcK+BkGZ4pdr2Odbl7skj8EUq
t4DGXd+2XbhB5Ixv9G+A0tIkRKVDChB+CETiWZRaNTPqBVpWVYKguDfUovoa7e1rBfZnimru3duA
L5h/L8nAkv/MwtS83PN2wjNVAmT6h5RlOHzlEHaig3zTPZ+Ot8Fu3oXLW7XiKo91s4PSTNyks0mT
wkQdFPsZUZr3SBrxLvF3NozeeUfV1r7c11xi49g0E2P1lHhyM0XKFFhuYmsO0uKficeZ7pt4Edni
ESIn1KNegUNOPhmPbbPuH8cOC2jgqD0eaEvjB+VwYlo15gKhFR6DRet4WM2WEUmUdcgyaoFof27G
UPaZNxRKMgKF+DzEjtazJb6Vw4bc2lPtKp1XY24WPxTfzrZwKSGejNhbyR0w7DpbBkepKM5oOApo
oNBwSDVYEVDOc9LD2hZ4oEpLCsnOLsnT7+8oNN+oBYBrB8GfHjLgrRajJkC6F9J+nEUAPMDxOQdk
AHfpbtwU/3BbaSaWoQmOe1K5KGWYk0wGOv69bdjvXjLrqNCjyHZD42XSnhPD1c9TD7aFUC7HEjHi
DABqyzWobqiwsDRYXHSApb4YH+2gXzn7NnK1OfPeMpJqRg9HB6ATFkuNjwa4NbFxcCuZjEfPGwcn
ANkJkt/zlIjd4U4hULjQ7aeNMrnd+r+R+XhQMFxKa3sfJFBSYOaLnbZv7RSO3gD3rUV3E2md4Oe5
IY0nuiAUrOBWPVd9IvJntW7OXL6vhgf9tvGOwsGyrucuQo1x3u/vLDYh0qsYBKoajjKz0e3ZH+Zo
1uGai+3OL30NmL0KQpI0zSx5gUECoha524mHN5wzHZZjYYOqcw85nLGNaPe6mGsQDR0k0uyVjHhI
Y4c56k9/zUhBY2UvzbDGHGG1g57Glldjp9f+AVnUG3syeZE1P+0tBaaGQcYWS3IvCiTPCWw8oGzV
RAjEI+cKTMWLHsReoCdz88yhW8mbQH0os11WgfeGHt22cUMNNvzJT3V5nbLvnt2lc9Joegkaop7V
MwXt2aT4Dv12h8QVgKcRcyOyEGCVK7cg63njrE5ABhBCxYRYey8Y55UpiiRJ3IpmRMwf7FzHpuGj
xrZNvlwkbaWOfQHpklWHq+pL6r+jtLhd/sVBeDDu4ZfnOrXdceV8u1L7ChIzngpkc7hQjNhH/BcU
UbT9F0/ur3qpeZ4Rt8y3iXYPTsL9HU3g1HvNcmqd9cI13zAA3+/Stap7kCtAhuxdxUSOlwKu3M6N
pYzleeM9EI+5u0L+zi3sAl/xQWBgIXAQR/m5P7+D3HVPsYwWywrqyNs+vkH9Z90alXHuPPR4MaTM
My4zdDY5sU3eb4lwAyu4rSmjWqWNSw95q0C14hS+vwBobef8eEdUGr22aJk40AGUkpF3n2V0TYxC
wOD+GoMAJ5iw8gSr1r39hrt32Fqf836Jka+B9upBUcx0gmfc3LEhIzxVWltb2v2L54s1OH+PeXHh
V3YELscVpIwcjdaG+Qq6w2CYKTPEtCIhIArbZcurteInfge1v7LJZljmfhGx5+wN2I9gjYpS5A7h
oGmh8yjx6FQ1UcEoZCv6R0cNv9htq9iGIwWSaZJLEbdNaP7zjDtXrDHrnV75sOYCczutG147kl+5
zuggcb/cOS17rBrRDuljTRIEG0nDM9oSolObPl6FvROhJgSBHiX1BATFn5QDiL6DsJ9pJGNxCz4O
musVefGUMCCXSQ+XCr4orGBYuxatKnO2ZFWG++iw4TnBPvdaRgg8uzvRJYbMAsFUFk7hh0En6oj1
qzk9S+JynqK+GITJhhIcaxp+dZdtmFeUvbQeTUR4IkKAfXHXMDdFXeg7qoEn03iP8r9Q8klrWF5a
3y+8jaNs0n3vSLiPaxkJZ3AmDgL3fQqizTIrHj9WctiqKEDKMHRZ3mzIaxDdsiiyn82oTwzqGFta
5XjSZyk7E145HjCKYb44hkv2vPGqw7QKpJddkXvHBFCfeb6E2TZyavt/UB53j4Y1jEFZbTEE5Hi0
t1HfBFhTQULpS700X2CwOMb5b8iHr3VdHkudEgzXyc0QU0Bi5HJOMPxS3YTlqXq+6mPKNcv0s/1e
1A07cn84x4yfia8dLzgUFzfyU5HCTXHAZtDb8Rk+A5Vmu8zkNMS8hPqIJ8qswA9EwVHcbDwkjOre
80o4fK3w1g59Jnra9vU4Wi1WPikneI0alt46YRRSfqA2EmsQBzX7LHyMJS9fl6ZZYOD9h2s8thjf
vsnvaXIdW3PuyqMIakrqetbFIZkrEDBayKmtG3aXNsq1bmHnks0lMW8yvOwD+pmJ6FWG3naGisBh
NxDvrS2LQd1Ul+9uU0Ua2taeKm9Tv1oHNspRD2qNmKXw6ila9Md6gCHQBx2gQ2GhuxI3kN2qrz4P
5rNlux1zNzJwJMTugDWdTbppN4FJ5mhi4gSRO27JHYT8Fq1ZmfcsqRTrRBJxTIH1cIbeRrHuDS9P
W60DMAZP5fT2kZrog1jktkU/jQzBH1oN56VSR/4Xev7M2G+1PFMs7Wlgl2gnH1jY3VpPBKJe87NH
NQ5RLyfEHh2WIvbmvebaIS1d+vvdsy1RYB2p9yQprKhT5zXejqN3zLBg+oRoY0uU7l0mIp+lYfVJ
llQwqLZQ5NUijFxCvVDa4zND+jqJZvuF9j8Y99WHQdxxwNssk4278+tfXwexpBamPqg5N/D8nVuF
/gISxzz7t9EgLxf8Go2f/JUloP1dOIg/UyLKIPaQIaYoW/svlg7rfQlJn+inIiYrkwUZNjbErYRv
65TfAjnnmWF/xsB9kokrhK4EWxIVOaaUp5lv0ZGAG4s7VDm9sLpWNgrpqqA8xCDyQJouB8hZMINS
GXCeK4DlKUp2Y0ftJjfG9l7hsE6rCOc6eSWJVAbsv6FQafrxpxwiocyUGT6IIup0Xv2N1LlHhS1f
gwbVmo8Y7BXTIJNdJi+IlRSHEBrzfcbJXja/omm3aN/GOSPek9F5bySVFkf176FxhQHpHW4SoIHz
1KtYql9LzEvhrenCfnvX0d6vj4YGUmwkYRFZX3XUkejvjTfYXnxfdvt8RZkREV7OxmcCsS92RUr1
sjzpJoZ7ZIr2FvCjE/q5DEJ0q16h5POSTjMeOciGuVefj4FkMkesDHPg2FrUV0xYWsm0LX8kAnF7
YX6XRDW9cgkp9eZ/2niJYctcQhfAKvVc87AaDUHuQ+/ZNrR79ANYu/6rErcZcf1MfuF+Qrl3NdmY
1q/KJGmjTCqcC5lAegNvbXjY7XYA1pHackNRjGgSejK0mY+bV2N0CrU13azgSfsHWask2hnr/pqo
7I9Sla4TfkjCIEbVpnbZNKGpA8V5w6+HghADlnt9VHyB2wTRyhcuxV5KuDvcFVzKY+rLcXqI7cnP
lNkNK841QWOxqsc8FcOpFsnWQqJukW6LPQy9HVSyNtwFnc7EMb4hTEJEvspcTiRCDBsW+NWaK/uQ
prWDuKjP/yaRLt+Rlyd801JUTnc6p9dOR2m8kzP2wrlsgcyAc5DmhhYbALwQv77hTyQPVLRe8sj3
PBUAbY17Y2de4p689t22jSTKV8xxRuP2/pSNEtD6Fdrumn86vs13SNiNMAi2UiKXiaEBnmPQUt+i
COI5nfN6gspbQnQsx6y5DXL9g5Jrd9ejYRjzQHk4PBRdBGiYJRPpB3ToNVqcO8yCbIIWaYKYXQRT
SxOjF8pQRCn9xbWJurDfKctjH/Ica8gdGMRPrHFmMtMeZLNXmgnGEne6s6JuDOcGSauuYsnT5G1z
byUIeXgRHgPFzFmptpNWYw+T6WgoMxRigucKFQyTHMSn5Pm9iOuP6kWsvB+p27vz1MCYRrM0lYl+
lLdH/Z9K6kdfbNdy6yKSIbE6DUEAoDx+L0C5/mszt5EtOjYKhw6OAvVheLw7u7L5r6tmIzqcyW3V
fGlJMY/x2+qaSH3ZoMKwJCzTQF80KQo0A0Idw8bDoEWrVIGvjgSDn/ob+vRjIgYSmAs8qBlxcHjn
ZFcF8fnUE505Hl3KdDuNjBxE4miuCVAp8HbFQNMqcHutcPzXXF8Llwdj8xxsmtvBCQ5s3oKVJftb
D1r7gFv8lrAIYKLdg+pTL2oQZ7PCjis6w69iGJn+kf2EUPGuV8eP6fqZ0qWVndVtEgYPDT1HCVSZ
2a4tAp4zu+UJ6G183X5zraxGUYt1i4RLoExEFOZLJAWL9Bu08HxXgfIR/8A6b9N4OinPFAAJO5SG
BPVk8Z5+43JIEB9id6UFdr2QFpjZuG9opMAc/ymSFbIEHBn/2wMhUNXJUGSerXh7ruSgwYimCYGy
9HxBVtrI8+BP36+NEpm8wykDIAjc0ggvtL6cvaigJuANfHPrcNT3Cv1MpOiEufDHHnI4UfSbtyRL
6muu4sJfS+Yv89jKccKcNgh866HRMjdRVkFQoUwGUKAGYHbPd208izlXV4EhI+dcZ4nzEJNKToeQ
enUMeQbRBbKhNawynRY5/smbwdsPzLeJDJbBdPAowRM3ydABR4Ai25GxB6BnAtip95G2JTkHko+x
SSacRMA+SZxuh5Q7t6Q2n73KhJIbiodetyjfttQgvOLpY2TSCYyp5PSEBbxZgKaWgwJRJ+sjGbbJ
fW+QkJmkXsuv4e8dweFJThFWFyitNH2MY2FJakD4C1U6KyzU+wPhb66V781lFsk2VueE/GD/9HJR
wpXDJDD0Qqp8FngAoEv9PtUdrGYWPnt6KOdOPuDRGqCVwTJ6/IcHWJk8br458G/fRfOXKjQ11/1a
UQ2iw3Elvbc+B3hR3MzdGsS0bZAL3Bs1m53OdxRmky8pVoONJXB93CMkVm9Wv0Z8OKhNNxW3HckE
FbDtOx09G/R8Pxhe1ewkq2Cq3+DFWHvQSsCm8W7/1K3aoOWvIOpzCsCNHQn5Ua39/J00f6pdld0g
sUMVAuQwMKeLzeCvHI6ZfNyGXB0pD5BB/jUPpD/ZhBHX2Q8OP6Htc+qNZhv/eEHWAFGmPF/w+vgB
vOeuQ6Sim0Ljtvs4Yy5hZhunKd4imiAeD+UmoHigBC36lBVXibC2LqUeePWblDOM/AuAFUEcv0hM
srpGNiiFOOTBGt54Pe066ruNb9ZQL/7mPYHqMzgP8ZROYRFBM2a+on6MIzaKes5ZMiPp23HdWCkw
QH9dJV9VxpgQndbW45CeFn81qYd7l1YNb5tlvv/yWe6g6V7vQmaBABEZBVZAp3K8RmJDp3Dko41M
YNGY4CtOIt0SgvWMm9xOS+YoYcq7OK15fVKMD8inCa1cPxRIJEti8YITbDB7B77QAYscpUJVbiRu
VFFskdg4IwtTUBpDj7lC0l1BZtQY5pFInRk/8bcvGOtny0rCGsP5SsF1N+9IgxyNB0hoIeTo0Y2h
WGjsKufc8q/u6Vmierc0V5M5irzfZzw9vl6IFw56eR8jsIp3qMsib7sA2xFdE4TkKmfHG6qgMhuL
WAteh1+I8rGGr7jQ9/xmvL+h8+L1MsnaO85yoExzy2fR0GwFYOXeCcnwD8ojdwPH+PTo0667XrDU
DFL7TcPV2CA3DXQf2bO1Ip/pFXdVZFzh29pFK8Q9+VB+9yHKBj7mmgl/RWVI1tR6ts36r6JjIBa6
iINGum5oGUCc6bohXlSJWmRCU0P9lVkXUM/jlCwxw/0GndNT/uo/C9m0JfEipLDqxTFMMKLUWu0u
Ochi1dkFisfQuFRyzMqEjNqaDBTEc7UXVZu7jptbiFbcdsTLRP3DV7zW6zDyVrRk4/cKv/n0NVFP
Q6j3ugfcampC+TgnV4Ge3B8l+hWjuChTJZKI2L42adtBHFRw68j21irzMO1UqwKafQBwETPvpmH4
TAuZP1aIV+rE8uZvnW3NNQ24/Yl1hqwNJJEkLiSZ63Bsi9+v4mY/sJ5pM8mIxeM1zAH7nZKu2N8u
ESERrni1LJLtb0DtFVhMdjYQycmWo5rBK9btkUFmQpqyYTQNuMDyOe5p3NdnLea8DjYi81Kuq6fL
xfI9d4pu++ZrRJOZxfvXEjmvvKeMn9h16S4/6KGNeKfNX5NWkhca8OLfRIUV3Sd/Ba9O7pZYlgTu
JxgIqCOUdCtlhls88MNO5Xn1cKM+4bhwkXIiWjPX1ugHk5RVxrWnRhJRtzxyOjsl0GTBH53Abe9w
JEoiIqWbBGjomIIfHyp2n+9v3R/9iDF3AGF4d68iFaRlRkptAduLP3Yr/VjSBKAOyowBqNMfqaIJ
NN80qf6HVTqKQjR+aVCDY5eutMowfoHF+4v4XdufFRkeaOXQ+mt3sGM1vCBbcmQvSJsF6sCrMrw+
MmWCKsSa9XPWDbGg5rJBD7Pl9kjJEccQGwLmNM64/QrtcqU1+mjogLwF80ay0XWoh39libQX/0Wm
KzRtRPTdXvWkHo8PO2jc7lr0gdUcHzHeEUYBWMBkdp/MbPRlIKc0ZYMHIGYK3hIg0ikJ2pm7EFDj
lFEeUtBHqocpbQUFDZvdjW3zgGr+4ElKj1haahzgwFF63nBs4+SahwgMaT3DgrW4/nglPT8jM8lk
dWqqqgInhIL/sqiZqDzPT+qcq73Zn1qonoIC3UZS64bBm228M5hjwAxnM1I3BKFURMx8js3WZ/2T
bMzIcrFYQd53eZ5avrZrTJ/NUD76z+q3r7oSiDL3br2Wd+LtCpDaz6H3l+/gb0wDvaWN0yFco2oJ
qnwY4p2JELNgGBiBkLJl+VEJAYZi35moPRYgHI93MibRvZNYfHNTs+QSKnWwmZ0aPpYgis0PUC8U
OTzc2QqnBGbrJYz3Ip53QuHUrhdYXVepASBDINj/VMygOuHvd5MNOMSupbPnmJmH8USLj1sqsenG
kr3uB9oUwYjCQJSlVcexwhaXSZ/spMyhbGd1kAq28Yy6deonCOYfkxG49WmkpuhHf9QZBCwHh9Vz
QcnrYI+SvUZzTpQYmmQT3tYC/LAIIDL2FCQ9SijAC646Zxdx9MKhF/N0uxsj9jmjWvQTh1uo818u
mG/gZx61FKkrlUOa8XlYTNLkO7cJm2JySw7Ao/HHA847/plMMbiJJyYAloKw9ve7cXqyvKWhaIvu
CsgmWzd0X+nuFQ/v8TI/JiQisBOy4LY7ZaJAY6uDwYESZr7hl9ztQ4Q6/EL+BNl/gxhdfVBMITlh
tQ/+Gsxp76hpsHUV0R2plGWvq3chpTKHfSNBlGSgULys15ElIVR1YKgNZnNTuUQ2f9zwCojthoR0
Yrq7hCCun8xKVeVYco7Bp0zj5Vl6HXiSM0j2YEOznklYcwRJ6VdsAUXfyzwS0kPyj2/37JmOJ9rN
JSiChnlwX4cS+Nljyz/crtjBSI04wKMWsL9Ry7te240dlgKRee4O2PyZZSiOcVgEaoQRwxkJjP6Q
/V3+H4Guj2S1tkA+0vPUyZqUdMRn36SBIKJdSNsWEX6phf9+FUA63kVuLc7npF4drj4LWa1FrFty
59kY4tj7cOEKNUtNI+TCl9ojYnWQ10TWyfP8o3fCzHqimQ7WUrk7EOXDvdpZnpIb3lHfTxxNKmAw
yHrfLfEGpc/XLdbjH0W31/JhbLUilud0MjD/z8crfVGn39hXsVNC+NslobXK0EiZ9lkS0fnx2+Qn
oZlXnzagyK7WvYwzA78cLI1NhrncYnwh9zV2mrGCac7m8TqXpXXy+tZZRpLfOlcvDt5AHQgLGxWL
ddEu5+JJftgk3auILIshRyvF8l28iKF2yISO3I3R+g+uzvprAj5azqETSu3r2waOyWgAdviHPdIO
Lk5ZNBQNXph60Kbq24memTa9S1ATmprRI6wRFanrUZVfLPWNXWL5rwMivrphEHzXodEgLW1nh7zc
Jp/Nr5T6OUd1ytbMpZrdQyugEqwg/64Zk8TN/iwv0hXQQo1r65lTyERwZ9Zzo9d6sje5NXBKJyVm
ntV2caROMRlbGL9fB0OTaxFBvLJljt2c/XBOqiDkehTJarAH+YOQ+q77DwhtKLvGPVSWoGqnwM+P
Pil8RmJOhdxWREJiSfvtmLrJkO3+yhWyPTNr1uSNapR/Ij7ShU59rTfNnCR3F4hyKfDG4UP+8wJD
gZYAtkr8Vl/sYBAKawR83fx0HjJ7ey6wezgcwFtQymi2C5oNiRuXAD7+1EyK0J2kR5nzL2k6Wyip
FI2N/JW1NHF9LoNUvt2uyhDp2RIIhGULZmNApnU5kpmOPPSoqFzdkPxtrAJqdcDKZ9ezRqNCp/MI
dG8HaOx8Avqhu0fNbSTKHT8i+1Hwa2+pN6rKoS0YbxIeGiKW26YULCeG/OI6AK1WeQUSZACyWQhi
Y1WJTzbiXCP4UbkrmuANSOY/pmtXiq5umi0utHksznMdsPopDKINKq/tNERzLv37N1gzLVUnijso
ecHQTM+K2LoX3ucE0/Hba+uIOzimNH+fIbJOvP3092mch0As7Qg84ckZHRnKUlB6qFNFV6GFWEDC
pX0znpme7g4eskG3JaFBbJNKbCbVfn3dWu0quwHys4j+D7Qph/xkYiC4C+MJ2vb3Uw87u+nPTnl3
qJzWk5hyWSVV6c0eGEh7KWBCCL4y0tMfA2+aFQF1KJf/OxJi/S5gj4ovtCQmdVjzvjlpmRZp1RO3
gJR8INFarJhP8EbtUe9kyKizjY9RmTY2WMYQcGtlu979YbdMw1MnQsI1qqItfr3wM4PRshmsoXOP
j7CoxhOJmq6vYEWBdzZim8mbGcP3WkLhtyUE2pCGBEzePCH4bP+5uexwk8jDmi0LpU0jAyd8x1m8
yG4soNFdP61VGfttbJ0KDEwcPb/9+/hh2+NjFXaDskfX9+Ug64VVW+nIx8JgPc3hG3f09VzN+rMo
lWRzV1TUxA4xbEK9XbC045DepRQUHEq1h0cLGh1dgra4E/NeqvQD0nzdCsdFWt+EXy8D9nsCKaAN
fh1YBH75jsh54C1UH8QzxFF9UNKIgnFnYkttrU+wrFOVkL1g+J5RNDKViA2SyXyZxctLBrwr+LLW
KEIeSTr1yBtqgHRkT4HA3ItRgRq1DwHD3y8lFPqgi9lOESOf7Bk5Z82Aa05A8nhDe9z+t+auEMHT
40HlN6xjikgWJ8En32eEubMkGvuGFVMPM9xjrn616e50uGOB8GV/MbIOv13qSD5FuOLb4kcbDGvB
2RLpbd+yFX8l3Ee4mYQOfwv83qEUKYUcUDsLz3RuTxgHc44Sz6s+snOb2jkghrko+ONcA2qsn+Jf
JyyD06MquJ5T8hebC0BMqPaSpoRre581mjWPjgeTVF/0fFTDNJSu1CmeVAtUB4BCB5qKznGZBzjQ
GSd8kmd5a06KwALwzD0uJ4dULEkLb+fFWr6oOmB8d31DKEAykEHKX6K9xb+sm++44EaK3rn8y5qO
Jo5F83YDkJ7rQND+DwN4rYbtyXzp4KKNBOH/H3aF1QpXZ+IN1zlhF5y4JBo6poR7P2H1zVUItr1P
AnBukkNO+TJiggMlx019LOIZUSlmBL/CWqZv2j1Ip5ukpf+M8qaoLHOFVXRIqIygiGS1vp3i/6kc
z9uA2GpcF3OH4fx1aOG0iVK7HAQZ35GcA70116Ir9u8CMAa+7gyjOur85/9mqBfvx0/sGMn1qsBP
YoZT05PAzcVaTcjRL4IO8uLNzYcKqIwWJsdfdVYFgiq6ZTKXXBxPjQoaJVeRmGzClRP1G6k9Us2P
jrmktCjFs0mcrgn9i+ZaP0JotkwIEv9LjsvfwW8dIWINEFqktxwo6yM+z82J6/h55cm4mbKZeCMT
o/kV5WrzcrEqdf6hR1ARkYyeN2AMBCDH1KWclQ0bGdb4qTwtirI9c5UGpx/T7ZJdEMjjBgmXmvpo
tC+0GyoJeo3TEwc2iEBI9qpiqaMKnKu7R0nfTwyDKaUZLHZ6QtdMDcAW0KnbVNiK1MSByuIAR4q2
UU12RQFEx5WP7e3sd4pSNGlf+CIQuO9N7dghmFZtJLG9l6g9mhpzcdkAWMBq+hbbDfMJ5E29cQuJ
nkTe9km252RQNSsTkaYzq4e4yR9ecGTplTFNnwv9cTgCn2E6nujYkVEd6eElz1Ekm3vMdwxdXPwM
flUwqmOnS4OSNqDwTedeyiSiMDkZcKi1FG5DajESooBscE9y6hCG0PN7AL5DrQDQ10KWp8422pIf
TKgelKABnWe4bOn4xybmGv0+f01fWxdDzxdy2wXJOEp9dJtUkUef1tfqD8wpqAHceFFMQ87e5Kkt
YdqQlewt6BPNiMHLgUgNcVHoW0CHDuXGGbvYrVUwe/wnOx8THPXV0NUpp1DD10byw6AZGwe4TlbX
OZgmrELOO+8y3xQG/78caYyt/LZB9figg3luzMd2nOEmNmpBDXA4KMzb+ZebMKD5z70Lvv9Pfut5
4fQ0j+LW0QE0ZKdjXF7h6BJAbnmHppQSIP8COFuvboT4sRPxf0Se150LFbWpv5JPd9bje9vtOrws
HNOwtEoGt9SUbZC6b5ktj7JASNLm6wM79TxbaYBc+rUdrIR+huaBmK1OqPuU+B85fL3rhzApanTW
7ehTSpabLT2RXkJFZzv4fzFM0ckd1WRkh0ulxblrOa8wDzgRebc7phCNIJ8Ka334F2XKopFRq/cI
zkNiPHmt8Fw25Fz27nzbjU/LR8SscqrprrC1PQj1dnek+KAbBMEBDlnF9S5USbI4q1K8Y7RSrony
Y2dLOeY2yd7OzREipSGDTEE2RAp+/9trQtbbU5/OpoH/1xN9dOGLENnceZdj53257XSEhTeY1R3o
mBtG0Klliq0rRB5eU+u2Sld+LuL2nHNj6Fbnlr0LjHoOvidz/7dAIBWky+xGnYep9QA98JoSvtX7
c65lsVpn4WFY08F3ax6jl3AcP47xpAaj/Rdrc7ZzveVfaigKDTLf6Jv8ZtVOofjPJmwCZQ2cGT7Y
W++FatbM456b70rE6Dhg6tFaEO4DdPhvjFuX7eEgoK4xnL3BcrJygcMfTfLmq6WTL+oY3F5vs0HX
ZatqKdaNrPYAE8quThZlFRSP0C3EyZaEkuH0aD6PMxpd2UGBl+SOZLR/WBDJ4zUe60ekK/bUX5BV
ryPESdpoHPf/Yh9aC/M1uY/LlpVgxdU5Yyp/UQnxb1TQJYhR1pSfzOwhP6RNTNDPsIDtN28Lnhy6
dXGhP3l0MCMdY+A9FKKJikCudxMyRGBD8UeHvghXRH0FZ2FEJPo0aPEs0Qoy2cEVcD3vECseWipr
3db8e7/R5u0Zb2ErnZvEzXEoQSSbJpjGiF/YqplgOzH+mx4aGhNNjZfQ9hhhacEmOx7SugmyPCoy
LiljaPwGtIuS3ZMAGC7nPUIfspgjmV+fwhkmheq0HRKJZb0EKA98fHOVUSJ5izZwP9AzJ01NcIqG
P4t66fWaKBtZmvlBTqK/skGhJI6F84/x2E6TnROoloasP4OygYiULnUOhVg2ZBXD4mGhbImblFi1
0u1C+vMI0fbr/nx1qB4cl9kvefD7pDBhmO0LOKvH6OvHlYIKFbLzrTpBZZFlBb7FrgmkUT9CQy92
8tKVPq67g5LW5zlJ+b18pFKaYH3vMEn91H/r8LHL5jIyR5mPmvDgEzbKxcsr/VETxYpzoaN/LbnS
/sdowA8nXMxS+Pft0F8FzHJSGQ4bajNIIv1/8G09UpepYVuGh6ReE54VHfj1175w5lSsqQjHzJmw
PWtVQSUZE/LzDIG9fAIwHIhmRK7vjiQyVWAyETs/qFPr9aWnMNDRRFVjhD/Vpe34N07G2fM/621i
BR+vQumAcIwuTD5koV65xON6y8iaULV+oJkAwVx5wyNp/6Lbst/g4uHR6Tqd0AfgTXaVRmbEjTYV
yfCu0XD5MZvTRZ/a7fWlocLdBctAErZ+GiZpT1QCJBfOJ+ALEdf4oa02bgQtvXPqv95aVskoSGIx
l7dtmQI/6z9AGnNrsDt8EO7RwyLUaUMTkcY3SrSmEX6h+DAKaFAXsz8TiugSitXeHWw+s+KkC1X5
dxlKhfxwOEFN/HJNF0wB2A7at2twT2Hzg53JK7sCUmlZJzKbmzJvpjyTWes80XhRVjc/OppdtCg/
8axpvLswjS/YJ9SsaDtxKdpGwgCLQZ4/RMZ+uNiSOryUAMZSrfA1EC++HZTIFDF9bSMsLxCYZmFx
JQghF8xGELXfVRTALnvM0MRFQ0MUvVX05gwCyNwm5JNIhZQVUWIlVXlmiNP6NyNSJEyXC2DNqD4l
iBv1VBVlQUOb9b3q/id1KuGRUy79U61FN5gQbw1jpIsgV21bHzKq4ZoJApUfUwMt+fq8MMMJpmdh
g4uFyznZfRhkiQq2CmrvidHSMp4xqG+LKLATduO5aeOZs+V9ZdcBM9g2pAIsfwoN/1hNEE2HPHTU
b6MBrWsWhuFsOeJ2zqWowz9wn7gLYGFsUO6WPja2Xi6Q1IBSl5xf/JEbZsoOop5jElS8NTYnnAQ+
xuRPf/paGE4sgrOGcHHhIet7WJcToXAKTkmUQDF7NBK4PuibBRxeJFMgHvJ3Rz24zOMx+i5XNfNT
nG70V/hodCc/j4k1OEGmXepQtMB9n2rsNgBBzaJrNGBS79afGQrvdzEmXHZvPynnx0CizNDFFGsR
UhqOBZq1m0dNV4qRpl021E90GJXJqevyetpCQQh/fPe5xYbUlD+Uf3NdTJMTuZP6TZi3Na/WDrVq
lvq9OMLCeq30qAO/UX5DiYPmMJP8hC6ip/5kXLQS814DixW16BZbrCkuz9ETOFMTWqSNwrBr4txT
AmBPpWZzQf82v/R6IuuXB/mYF5y4XznWB8Xf4i2+2Jpn8VksiCw3dvqUoroXRpT9mxB5X7EvkQ+l
YW1WQkM87ig2pqLgTzlXsp0zYBAullBt9McCYgoP67niG+8Cbgcgl1iW/sQD+T1wfkroQDv6tIas
ZlsdgEwSXZvB7Th7SNi+5hUy1nSw5bssQrTxqqhTeIgsZfHvi4egF2Fc37Xs1mJKOM2BaHcp5xOW
WFWlNWfJ3b3Y+dcaCiZ9JvgZFJJXWyGZdGh0KL7gPPE9da74TTnn4EC3l8n5hd+OJ28cZfIpVj1O
5yDIJRkIR8CBsMv0I0xDgF4IRBD5OntRkMyVJ9zDG8O1yCQs66N0qbdhQ3ptEIREIssGIlUZtqK7
jfbyydOUdHaIZI9rRWNYoNWml8XJTKRKNt/XlKZN7hAVw8J3zoJm8G2EPnjfgWwIFvhpBNtc/QDd
1tbOK1Cd93u7buGexlCPD/R7Y4YCLTzTab3ioRBimKvorTJaA79W42cXvc/m8HNac6lW2zaCZewB
9bhD8rIRPQCfzKRB7Kd5d0FYo7DA6A8mhjP0bXFUP/uONGWhUbACLKBw0/Sk197HMG2agte9UamF
W4JPIQE0jnRjaUwFTkfIz6OD61D9LxY+AxF8COrRDlvEpAgoYEALXZMybqheJzmCOqs3ZkW/tW+i
EFLMEZsmtWT2py3b2XYbXMlci3fEv2JGLhzQI0E8qekvY9rm5NGC18Pxyz73D98aMWMBBpLdWOrP
50m4izWM808L4k/aFEZ/DQi6lKpB6IK4XtYc75qsamajlJfBW0/9YBvVeZSndTAU5TMRy2kTiyXD
hvSnevFKJs1OwuGgJzEcHraStK9hDCEDGAgNF7GtJS3EdDkuOYD0d9V7u/5ImFMtfGQ2xOX9sm1S
be5lOcUUp3Z1NgUJ0PjltftsNG14YZhPbpP1OKweEmTPg6wzIY8U9ueH5QQQMLhI2uYAu8GUvLUH
Q8aRsC6QWPRa40Elk9lhHIWrQJ6W0FGp9PQXoPzGn+hOZu0QzC1jOVsjeM4v50vVapmZxQETLRWE
/1OsBw3L37md5McZd2sMZTBVeu+nepGnaOEf0pFnl/dSiDGYF6KPuqnr6y/4YPAMER6J7v9nJW5V
rumH8zGrY9y5pc0F3SVGwBFOZlO/SNeRBf/JDsq/YPk/AYoJmCw0zXMRYLXVy6ZDnsD0MPDZLUAA
0MzhyMtxFsV43QX2ZdehtSDyG2hPwoS8InBT6Rq5yWxt+7RO64Hxyri3MYIal9y2SYy0ml3ZpFT0
9wwE5bYf8DbaKDNa9zDbAwQBPr7f7ET6XpKKV6pP4laDigMgdm8sPd02iZAyTUUmbUPNO5FeGsBk
pva5x1Ny83bYskoOlyvkE5NnRGZLAHpqHgau0j6i+gI1vO/u0ejIt+H3ydxU/NSMFKZM1NL7XIbh
PL33Xq3hn1UhaVVGD1OqHCNg9t3MM77yt60H6TEAZ6zR60jupRT4luV0jEvcNJQvwrPHoldr+ZJx
Vl/jL5oQucv6ovLpxLl6iEPdW9sH9swB8w7KuLuQXEU3N1x5gZAJ+a+m8f3w6rh6RLq26/23vpWl
5Pd6zXrrxyC8iF3u+QG+u9WvmSIPGgx/gIEpLxvO3LaXZbIBTwjv2bAhaWAsXGuFc6+fOnwnOgTe
jjv+WsmZbct37Yg3FKNteaMqiKVdklcsvB1n9V0XC4DlIMXNE+ZhOfyFrx3T5ZFZ/Ef+tGvq7Npk
YUjSlKBCrSa8insZethQLiKr4yRG245kycn5IaWywrT/KkTty1B/YgbvltKcEWKUrMYdE3bMW4WK
oVZ9qzZmHVM1Xw5QgxJ2Ww+SwTsl/2ZzEUTMariK7QMaE3CFHNQnz4R+6GgqSDAdFeJ/wCtNzBGr
fLPMmecwFSMJbkuaOelkm2jSIbEjFTreJ90CWoTfF2lgoKgzt0GvKwxP9Uxv1uBNImVOB39jmaPS
4RvDUuT795jwBqd5kiLGMcABXvgvm+oePvt9cMNFze1ibYeNcXioqrFd0r84KIlcQjOfcsQi1s8Y
0PAkPtkIFAUnO58MgXmaELrCLEbH1R8tjpe5RkHyYWYyaulD6qp26+UNovzsZ0bcAtqreRpB++4m
Nhr/oCExFeAutgmOOCmFANYbCh2O2LAekz50is3q/4HjrXkZcw2iGkVJ8zmwJh+d6V+5hLNnwiaO
vHltIV6OzfdcOtwhHlb5RJLbcyg5LXqKwcTiwSlGWuhJEtVul4Tlc7t0CbJgsMOg5ZkRT62BVYRn
EHChicA4pEoWHELSJ/w3tqGkaw6TsHFNWT4AAj9Ep7ZynseJb7C0+7iDnSMPRAMchuJgPaE5RJFz
qSiFjLPaLzkA5BdLz9HHINPUdxSMtPkT04gXPZrRLDnU29GkTqWEkdRFM2Zh01TACWFARq3TscxR
vz06l2Sjka/mmrh/RvHUcwiQryFtxusITIKwv7t1RmBgRpmDpv+JsxU5iRs4qe/klOsYz81RI4mr
FCnsZw4atqNvg0h90ib6Cd2WqsZwlR+jyAowo1faUP5A4hKKNvjiIm5UcEv9/oPEgBs7AMl9ob+7
OADJj7JwgeEiym9VqiCoLbPt1ZgnPt7wkPvbOkvtaVxaz7Fj43SFQnudzya98+JTwpQwMOvpVbTD
pb6cDNY1MIPi7NiBUNm2KbuFyeMCWsW2QWkCco2GnC5lc/piwaDSsGn9A+mKvliVNknHxG8qp6VO
m3eQKHDxsBt45I1jn1/4A4u6K98rJg/OkEp0AxMsaDyktK2mkCpVOfhUQv24AtZMHmwBqJ4wstWl
e0Q1kIu0X3R8zo6FJjGA7Ee/CDmFCq6zNgNWrQWtJeLvXdqb/tgChuRc14Mizxmk5JOCylJcEM5c
iiJv3yO0Bu75JBXSpMjFjgRFSYwVFLXbjmWkFRld78+/cPEUkEH/EArpSBlcVI3BYK1ADS1PmHDf
HaPUvNXqWtjtPJEgKUdUhjx9TrKAdn4VxlLPIixa0sZRL0QCKUYtiUJpALLMmdrYFSUkcvnikAi4
R8xFsApu/wgyKoa+nWI4N8fwgsd66oEeYqm5YbuvXxkxxbV3NoKF3nfylLZTLUpjfjjnlFGNFhZB
3E03hyxadgqieY1Vxt5WZGodtxXHyqpryqJ1hpNWcbdcpAM4PaGL5CYR3NtNxzy0XbPxVEeL3fYI
jhmOD4gHwAQ99Pb7uU+nYcoky8k5F5XMCBAhzh4nD/77BE3I5l1vkjgwiMqlXzoKRnUnUxKsLHBQ
svrBtjcHrOLI4yg3N0dLstdDG3OHh/V3s/AjGyOxYF6v6goZfBkhLaa7AMasOJemXRzsvRrIjFmB
q4G2OQ23B6nymWJ/CSFfYIwGGsfjtgroAeyv89b/GFadfuvB3xyib/nJY1URLs38yLzCC0xJ9gD7
iluOnlTThLc7iByJvGqjMnt0izZETvbQeOZs0ynd4hboCm5kIdjVhq0CDROn+yWdhrEYmU4jwGXR
VP/RaPkXXC7XDoJ5s0q/6JxkRQrZCp9q1ePIhLU97FkrfEgjXbUggoey+M+Y96adQPjkSWDQ8JAz
+VuZmr1ZZ5kNuJFZL4G2F73rp8cKDuQQfTuESUdGanu+ctUGdHNO+nNFIsIsdt2awc7Oc5wjHy/+
cTVR285Ze8d5fT0UpxPBSRLiFi3mexghTtEJKxfzBNBuBqKfgI47PMvSLmBuLmMJkUG6srDJmGd+
PpTkqbztBdO2nHiSAPpiC2Tkd6XaMXWVX6zR/NhJG+XtVjoUbY0nPtu8K8VQJI/k+DNabc15w9f8
oXsNFi0dGPC8SlMVHQR4ZiGlQvp94EDNgedfEt0HVB1N/sSac0AR0703HEY/f4k2YPtIopbd48WR
BBSVvWgy1w41su98fPibDUxyABAGNjeWd8ZCaPi4m9M1VeduR8gAabI5Qht3T5nfETH9dICDMLw/
HHyxjYOGEr9reqKFbJHsg8YURu2FI+ESjj0t2ko7zYPbkeKwTj2e1jxar7dil8PX3fC2eMy1IagX
mfVKlG6V24aNzrHEPi+yxlGUUwLD5Q0IONkXJTIu/zPh6mGWm3vTjx/l+0rFMuaR2Qz/1YZKz15X
7B/14cdDUf59liVkgxaRpte8GuBSkPnYJET0hDatLzOvycwwS3oAMrFnOA4/VURnlR5GagDlaRPk
b0qUCSfskaaM0HiaP23CY+SbwG9kfRTfTrASAQMaVW2xHH+gzZAyhgKSPFrcIDocWAlx7mz9mMor
+fotIVI9lpUL6KieZUkOfJzlsGGykDLn8Z4ZNlh8OjyIBnxUl7iYj6zK6eDzncuNKzgPtJBhBCM+
rO1TkYV6MfuxLzUAR36Tf15e97BRZ0JeVAktdieHe87q2OVaGbysFX0Sc5hlsivfcgX+1eoJHceM
zqHm3tL5Ou62nP3y9ikD2zO6NJMXW2n2t+K02t08jEWWH4xX53l1m6ZqrRcqfM+1f1DAKweX+Te7
CWKc6W48lUaZ96nRg03MzOX+oD/uNKvvgjGBD4f6pNpQyFI8a1smHRH9KKfWbJSNG0/pXun7z0dc
AKnZx5Y997gzgMaQGifk7yVFfHopj3gptEiA+ISf/I38zNGPQOwjzGz4S9d2TQrcQT0iU3UMpWjT
Qnzd1mM2KtD/16gHT9L4Kyxe4uoV9tsNBDOwWg1Il0k8JPw6ug2baCwt3m/WQNvKx7/Qbsoh0bhL
g5yjmHkUbMhmzX8RZgBPSdMeKNuj3sxMWLLPy7Blm7mhEnQLp5Ch9Wop4fL9WNDlYEAxGScwCeZU
brfVRayE4TOb1rn3SpCRmrZdnjoZ8RnX0TrCdJKcxfkuDs/VZnB5FCj3K/nUh2+QH0zUeJ85tX7r
jMDqkSdt9hiHlkU1ET9fUjd0n5b0ojV16qDGmPAJdj3pC+Br9u1h4XX2uj1/j+YIIFrG0dnaiib8
UGEqTavWxy4YDcV002Pz0ddyxjWgRDYfJtZj4mAFZ6NtiwfAerVc2Cw4s7+u6fT/doz4onUSrFW8
HhJZY1JOsLYLBnD5dC/xwzpiWas3G4/iJHp5lEPSRB4pWXbYCeCSIYN2jEopdzyEnWQOmqsg+U/2
IWHWZ/Q7dP5KP9R6BKLY2ZpLdnfiXi+UOxPdtPNdRApz6vdBD9/YYbqfcBoLByq0lEqJn4++5pHd
rKjPCladqt34RWHvs4RBIKkOPFrlZmFlXcbkz1wD19r73dM4M6tiR81LG0a6eMpxM0QwjcG5MyNP
nTAOlHJmsAHuwQ//i5OiLxKTjFA+T4TiL4QYYqSz34/bA7n9FISoV4oekWXw+DDBfl4C2KXplAPW
Noy01r6XCDvtZMImfyYuJAQ7vxKgsTgaWo0TqaL/dFCM1uxhvvOZRTfJD12tO/pL60flnzltEyYK
Nnz4DKZpoVVryDKA4sjv8fLWuT068ebUYuGs2ZqAU/RP9TR31hj1N0N5FAR40L5gAv+pI9H2N6CK
3jzoM+p1p4ZNwQUoAonzBaQhmw86HT70VXaLqwO/aava80UTtFSx6gw3iKjvQb3C0biE1JcxB2G/
YBoMI5voedVPLXYLUqyUcPjRuQ/wGnz6He4GgubVN9I2g1LyYjfBoc0VZjUkGfyInlmyOVsQYP2i
z8fwi0JV8lWIbnXAynXwzJ8+jZMaPmLNjc3ikSeCtGXSsA+rJw+jvNLKXiMemRREIuYCPmA6bGnm
fNjeloCIbnpXZK60lboo6Rm6ClRuzeKCKM9nX6sZtuWIfyTIwGQeGykGnieMg4ZQc3JP8EJfL1Uv
6y7uB+SDwNSVowBYPkdnxiw10tRkooNSiGfgI+Cvxu/7pbk/tAJvC58OQpCemDpu1hogkms1UPqg
bIukd2hFxru8+kU+xvpasZA3EFnWPhmyuYl50YeGV3QMlJDFu61tbYyq8L+lMtQ+b9h6Qr/W4Yfy
E0kw2aa3mlH04/LgFzF+YRiAlBGilY/Qu7wdJdbAkKxrpO6i3E1ixQhJKSIAv9V+FidDTEqYorB7
9zqZY3PB7PBJY9YQ8+qnrmX+T+9VJcF90XsKkUMsxXG4cT6hSrRPw8iugMflJolreGqhPT+ROigT
H7U2A2wVhb0SHJk6/C+XBanEcOvI0fphtfOBO/JhW2kvn9R06doEiGhNUe7ri4721KUSYztJEUvr
m2RfV6Xdc7Cj/WvQiqYXwQoniqNCku3cCeKrUuYfvsfTAoV2UL4LWGUuFriZR+FkkwKwI0Vw5cDU
dlZhMfWB/T3jFut3tadjK142iUdFyTvTN6YAVqX3F89SzOLo2CEXXPvdB3r9MxUprgJhSLHx2cUf
/Kgj5PJWwnEigDIdHdzw1iunP+ikp+vXNgQFuaABrILjHuWcMOeos9LyNXe1TwUHQnOGlST6wjbR
VPqxyf8OOjaCAgYEFW5Dw6r2TAo4IsoosM/nUqAutSC2HoayyBkdpEjHy/8uZakLUWu8AUkokvjl
w1zcb1n+aVU42j46+7IEhUWbdA3NfavQC/lBgcGuZIx400L2YYG0Q69P12niIypnl+3YLlf6ughZ
3cVsZ+hpM6MlSSGLLAoH1qGL2i0950h8U7BSqPuC/QOnFXJFcCceKoHYeZnz+ugwFxGb9YQundRT
gQv///evrlTAVldkC2zPUju3GPShxRRmGrinmMepM4HSPbsuhy3+KwCwMQGrcJTXjGiIg2oaMv6L
dgIiDPYdCEBiWdnkuh8oErNLlXZHZGt9u2MDtTHrDxSX8TqTxmMeRbHVhaE/mMeFKhwViZIPTWnK
nzYcyt0yR4yjyjnCthjwHSTW8mBzN3TG/MQb5GfOyW+DPAkqUjYKZj615yEBaNKPBvSwQxWE0KwK
LFgVyortqfSLlfp1D1kd/GKIHroWxO7mRNdSYhdVxbyBCReGKd9UdUDwnKg9tw355bdklq0RgCMd
MZt44QHJdrbWts8HB597H1jpUvA4mEhE3dYo9M4vFcIPFCsrCIfWn3b1IY73KPJQDFhiwB35KoRo
4LF1NXZD4+/4MUCMNaMXnA6aSir0MdG7zYZtBYtaawlY7mkBVOCGAP+/Oo6uHchJ0ecKu6ptgeax
FkjeHSjgyXs2Sye03o/eIv4CzBmaaVUOTEaKk8W+wTevBA7dzlbFOvd/2e6z+1YBxfdO6YKREKld
lZhGZk+SyY1sKoVpfwG2z6I9dbACCKArfGT92z//f+Wnsk/0F10tlq3afM8yPpFHxXnVIfIotEu9
V26iyq5UnssbecYznD3ttimKrsQJx/PuHALiVrYTGKLPa2Sw/Tvarcx+lPBQxt98WOrzvqr5g1p3
Zkb8MamcfxfrBuxz0OCF+PwtuhBtvOdz4ylKeXr2TxUa+pHU6qTV3JneCt7+jBHRDh0S+gS9445R
CWp/tP7PUNngmwNdVje/Ad+Qwg96evqQm4F38czYtzllzBk6jfIpMQlZ9250PWigT5ckJ+sz7OeS
ojgFHceFScFNrvfvP4FcjICMxp+EVbT4pLf9tkIBQYuT3ND6aCPCspxAIK6DQpquGDnrjRsJDskJ
uuYoalZiLr/CtGl6FAN5dWx7Q05gqwjpSrhSLubb0xCdz4J8MhUOJlTyvTV8JqgLBZB0hEddHJyk
5Huieyh4+0uWLFAE9RR23VR1lZbwznDK7zlf9r3mcb/pgYpnrqtIrGDfIq9RaLX/VwnS2wHoztEf
gvDX1YkfX15JJbHEZXQomiL1u0ifk5rjwiJwbwBIeyhuAlj+nHm6ObeMjlwmmDODnwrNoBLmh2xw
iXYABuljrlhWgdCIdmk5j4DzYLL3EFkSOdTOWLEn423Cx8/OTPKC0pM91V4DLu50cyrtNo3BweXX
Ey8t6cHMVeGt+2nFRaAaUWz1oL8qAlxS/I56X9IyLXFg3RIq4+Y86tyk/0Gtu5EBm9nWQNL+KDA7
FYwxhoEwhGwd7iF9UkfEZcg1GBASXKl/FN9A9WCqe+acgrwIms5qykJIDO081/9qximQ7rO7doUP
uTCH+qFcjGIb86v0SRgKYQ3t654TK4fpJZpWK7PlvKyyEQmA8KE3EHpk2Oah2ktJ6GnF3Zdn0vkf
uaK0hW9IbUurTmB2HyiHmGgxuqarrlQfEFZt0aFWsfqPp8ejD13C1IiXEGG+8oHooYOciv/EAcfA
v+1m+45rE0zKdxpbugoOPVy6rsXL8SFf57zl4GiUiaDwGspEivr/d87kI6++EfMG4/2EnV1B0kp3
pQYnvaY3BxnJ4ybX96Jd/QxJ2DW6GaQplrZSl0i+pn1ASqZ7BL9hs7nV7IuSKhV70TbZI2fqEpeS
4oZKsBz2tSd+AtuhufR1al4OECaSir4X9xjsDIFwUEx3KvVAfPB3zjxzklBXJcbdwQwcahgG5j+R
QZEf1kaBLzpLO/mVTN+2wQ+iRElvm401gzXb5T3trZkgEqr/a8FSHrX+Uy9Hmr2t7b15yWtNrg6S
6JlBsoJuPRMQNBpS9uEcBm/D515s1bwxVUi4zjCDbkd5pG/1Y2VWuoiz7j61nuuZVTxC6MGXfgEN
TfkYrzdcrqSsWiXhlJY+NPK3iMTDJBh2RqSDcBpMaWUB//2ImXznLi8TcnNJKuilWa5w6ux1qWos
8UFu0M1xRRMVd3Pd1n7x3jvWlE5qYL4jrPblTTMGEtaTIdM9mw5eRRd2v+fXsGaEzqaJBqcJ6Ahy
lyoMN1mCEN02pMRRmJBkicHTymGPUkEpEfq5AfVh/qaPBhnWY9JdJQaG4Mq3Td9PzSsakndtFSxl
mvUqh0CfvL0GRKYqapI1cSoZxtwJ7QgaXZotqR6R8WyF1vCkFSzKdaM4ro8GZzbAkgkE6N1cF3Xa
FgGXIzJN3Rf211Eu8PtAXN5RFMQT8AFDxNFVtKN+Cx8YCP6Z+vpNh20HzRuog6SgUy6A/aBSNiEy
XRPA9HwrTVRW6oCwIgLP4oCPomwnKJ2bly72OILqS5UlVgJ4beg3C28YkIbO1bHenUSReY8t1ze4
WD2cpOdhxIjaj5pl34rD5xOd9jDbzbXBrsB28UEJM7+cAai+16uxvCGMCLpcP8lvtECr+Zdy38Ds
iFhyWN+sFfnA5Hc1/XohVZ5FVH95uh0mVTANMpiM0vEgTS/DjRIt1r+ohvHieq50MgLrOmA1GW9k
KBlL6uLQF6GK1DH8FjMTZ99OvL3W6EFTu6vVaYSF/OkHi/aiT8ZVD5QYsxzQz3tDrft8C0X71Km7
Z6QPlTYeYqblUK4GvE+1P6V0JJAmjfQ2Ix9tjmv1OhHyscQxdVmZJdcAzwuMjCDf7inBDQdhGChF
TI5cn91RfnZKjP/77mxWC/vtKXi0h0w5H7Mwxv1KNjFoEjrtuuT/8LadK4Xdva7S766eJaCREoOh
7mHZJWyb4sdZCllEiZT+WcxeskCH0eZHXkLsxfwpPS9qHlH2gtKD3BfSOrUM6CjR3VS7mswdZmdx
Jyn6IYv0eQc2jJlA+o9boBcMpO6AJybMRouqM1VhMYPp7STfmyjbL7Xl18IvQPkslBz+rksqlmV2
/3UeHmwXGbrXhfA/pcgEidtGHo95Dgy6aCrJt4F8tZl+qkL5LJwgtM5ADBuF9grRua9EClwQuNyN
f8NpLk0QeVvpEa3aBTAYET++Q35iPfx1oSaszCDaNCHG/KnXOkUSpPDqHmPC9ya0Cs01h31y4xCc
F4lO+3gg9MK7iLHoWWRs6GeI4kr2PY3yfApeHMorLfa9DQOvOGrRmRQmk1vm6HvqsICR8lchdcp7
zGQhRx42cMC3I7DxxAlgkea+kd3Kk2lTuEexsMTt+e9E1H4uCRtcei0ndgbQ2uQcgUlo2IwxPa1Z
OJk44hVHj/rIvtr/Qsox7beJZedMDqLRDofWvK2KYe8YBRJX1R1Z2ZVSQtvJzrz3KqYj7w5vzgCz
1v4RynZogS9zML8RgDHSNNkKcOn35Z2WoAt2+r178SPxL6yGw7vTq5ReJcuOOKzob72/3hPXuPiO
qX5ZAV0NH78mtH+eAXnT+/W0kQ9LM7P+a1kRhINtKxx6MUG4cno8IUiqR6wt0qbnbe+YTKNjvQRV
1N/w6BwA8FSxTw48RJNYQWjgPky15jeaPIOYBvpBrOriCzPqtu/SC9P+Nuil0TzDeDAJROgCkgsh
lnoM4OtWTGbV30vNJp+6aRD3rhDMgWmun0hqSn8K8/qq4g550jZKPlelGO84WzkjTuSHkxTWz9v7
DMu/g3qExlV7Y/iqZ+81g/l4QOy+/EZb0K0BY9hGpyKRTDy7uYcojRToPI36nK70VU2vrRoPGK1o
YITmBMfA95RWpAfJuwEbWBHQknjN5DuO8WmwAaAmA+WQzYdXYIt+5f0D9uyfVh0MPCXM7EkAwsSM
sZo5+5Aromiuqd3eRrfeF2qVLX9uO+iDBMW5Qn/pEI3AE1kTyVUGi+YiGTvWVHm3JDfzC3hfO206
CMhBdnzd2LiElzdh4SVRGARN3XITflJ8U/zzMTjCqUXXcbJoCHMNN+gsm1TRWs23zXMbFkNJCCpU
xQTPY7Vv7rW3KaET8Or7lc68vGvAZV7cr2sdurzKC4wyont1RhnzTvalPLGg9Y25Ugs/OU78DABz
WOaH1y0MNEt/oV+uP8ehTN8LIY8wN3piukGTq9ian0xtRCGp7wkeBO2ivtFE/WX9MMLNlrPHrKcr
ZWLIbk25VyV8nm9h8bYNFTNTwkq4d2t+9TrStol8OgKeyrEraf0u4ySJRJT5I3H7unu28L8sIbTx
Y6Fm5mEcS8PbztVqLiCS57jXKJUVq2AsbK9cv4n1Qsypt1ER4HQBaPEXnTv88bqcNy+OzlhVgQCI
fUa5e2VUWYEM26rKBKamLSRL31iMpBnr1RHpiuqwohoGGXR3odQr6KzTNvuajYH/aPquadZdcauy
RkdApe1tPUdH2gSGHYlcXyXccD1B1ekn6JND0r+SB++AM2F0KBq9fmtR24+w9PJDLy97SZYSD3z+
I1kQePrTL3Y88rmSEYWPXxxjeKrFE0UdMH3SB0acs2OQqp3X7oHHEYzMIF3guo7mG2Tf9MzVge5V
K6PDA1ctebIgwMEsa4RIw7lzraOgSsJHxK+/Sp1X3VnRVsqggsI/ZP2in3TXuUgfpg62+eh6bAUN
iVmCSZt5hW9QTKOc3jX6zha3B+3vK+np5EjV3DVkQcOwWQ7A0au65Li+EjyDd4u7WhO8/AMFxi1v
aA3mYH4GiRqAwqszyBub90TRZ1/AGTnaP+4GrtYLj3mZ+sxJKPgIV8qyjDFUBcCR8IVbHulXeYpb
Tov71KXmTkDl9x6GHssq/0JOs7U96suaiXDEOY0R9kw6gzpyLEVHRuINl9JzuZl74f1Nx24JCdXB
QOSRIUr3Uk5YrEUdYZ1k3C4jhBgfmq4xz8/v490XtASlL3kICoqYo4uIFZbhh3WNvrYVdqckD/tj
qgVTtqUG7GgFiKe1vpF1Sd9SjhA4NlouhOSQpNEB2bOFVW2qSOHtDdqMFCnR7P0cKTjFd/MYewFJ
JJFS+kZCQKM2TvgvR8GY0CIN1FklIzfkQIh/2v3JbR2j1zt+8tNbO+L58ByQgZHXst7ZKudbLJGV
6DeZ55AkJWFzOtXGW5sboMr3ABZwB2ZhbwpTTVcotQf0ALgpeMmUGzxy6wzHT2Jr38oW+SZJ3thB
YOuNXnPHC5NcpyVkom8iy49BCaB7cjZ9S0XCvcngjaVbxq/7H81/KTpCra/tLx3LxB5gtLU6jVqi
VgCtKRnymJdimWGZZ+AQMmpi0mgB2Hv08x+asE2nI/zYp4QWn/yLt+wZ/zhmomDNlJcz2oVcmCZc
AANoiUp7EDVB67MHoGTrJtbuXsqBvbCM/GwUNO/Oxom1War2Vwfsrvc0+mLYic05qC3GuN/s/SE/
LWKDqNlcRjb8Cm6PyAD51v3JOsLx5a+aPv6NX5snxBxl7Zay6OFQFzUHHK+UWA0fPmSVOXxXtUPz
FODaeIzRgF9HTN9dcsrBbVVV8XlGc6eZeA/FKKh3x2qsZ4LFgmnS50qGEULXlllUveQhUhn81RqF
kK+AQI4D2kZqLonOJHgCRclJd1NjV1I8Ty8d6J04oSYY3vDpfOWcVlvIOqxFX9VjyRya444i0Xp9
jntF17TIIWP0wOB/WtSe3fbYv67h+bIAIosouVieWYzcuMc2vFYy6E+3H9ju/+cn1pg92KN1VcEh
ZugK7ocf8o+TXz7g0m27XNds5oeL5wsGQZZmD8dZt2RqNsDkEzjvKWqA0Vxouoh8H/5c3g0wWVrF
iV6NCaSU6qpAH9yUIb/s0GTgaNbdPQDHgrwF7jtNC1y78FSF8vVseK+uWPI93H9CGJVaYKiVJD3D
WBFU1RhJrawASjIQTUngR3Eg+MSCxA6R40yk0t1i7PA+a2aqOmTeop54Q+38LUOJywQEj0WbJjEB
0sutzSyjoM5+G/V/Nwp+G+EbxAUQ1T8wzB/UnnMP8inOsHEkePrGklcNGWqf9mvyW8Xf+jkPWE3f
v06rXGIwHqQSj+C+AYx+Fq4OK8Hki5bS6/auoJU67Q25Q5/3MJYWCWbKh3RIV570GUvPpAHD58Wm
YBnVw8wQzAptQDh6fULxzn0WMo9iAR7Pq8BzFh78S2AFvhmGsSO9bTlLlx0JxnUKIbT1xeBYIQlW
MqT/8rXDEjfMAQ1cSYKYm30mkoMjlpCINe42rRQ8dnKibkDMOG9N66W5A6VfoQVYsg8dlIMAR1BK
iyJe+y5cC9yAl0LmbOygrf4GS35CAApvTeN+JZuyX4rG+TaaZc75SAmvllWuwnRtfakStG2aJ9qn
OyfiuP24wXDLEA5rdlFUY7m6XhYcjmccOwVjicupy2AOFpn7tiYGhDWBCmSnNBvDPAoWi3o3/1Te
gVC1FALDkb6SCHyL/mlr1w9CAbfJcFEs6VjZZjR0KRGSAuh0yDhp7w048rDZWZBaAJfrtZe3poF9
N6Vtq9zhMoIYDhAARKY4O+3o5rTkwA3aBgBMWGy81desIMDGCiY5H7e/B8mRoAdTCXcq/VOc7lFO
4NJjh+jogBl4OH8m1sEvTlB/OWtqmtB0gGGuMdxqNRkfHMR1kzEyZVT0E9B8MNYf8uwJNmxAeIyz
5H4quWTqPk3qAsNsW/x9taPiXxJ0+lOYy6c7SRDeifvD97YaJmw22J+iQgBgTnwQrRszv5RDbVYI
tprpcc6oz265ITqSyPK3wyVXDyXeT/e1e+dZrx4bdXbViHRAMc0cg3dHJ/oxsi09CVi7B528jev/
J/DmSxqmqOYb8Iq372fdnO9HVCUJ3r6chuf9pW1THifoY7PdycbyTlXv+PVnjSlH74tcc+4LnQFO
1IxsjfChDMOGjNf9htVpQ8mi56WZqo5Q8pGQ1qFxqM6c0R4NkSL5OhCtWp3GfgrcQbyG7yb/W4Vd
MplRt8QCk2TULKBp4oNxXpuVMvMf98Fl18uBUOCM/lpPIbPW+kqD3ocgRNZ3CBORAILCcF9fIRr1
t7T9zk7MEzFhk1x9BPZpjNXGNADQ3E/VK4wUaaHXIiOWKSCGAlanFtfakls6eA2NlTFl7gmmy+EA
+Y9rGV9PKRiOjX64Mbxcu8Hkwz+jdg8P2QxKtarqJcTsn4cWNj1JDY6nYKCtS4zMPihIuLxMbGOK
PPT9HWkHNbBpFcKYvk/kFfL63jtI6Ddsw2R1nfUTjno2HxTNejidqWG48um8zaz+ujzOijgUxVu6
d4Cr7rwtMZmi7wgmIwj8k3SQ3srL8fznegr/VLy/04LKFJZqZMPoanzhCTa3WDntNBuUAr5dmiRT
PHXzixLpXMPiF4HRgaWRe7HNLlHc2IpAJa6tVaNQ+P0lLzpfmDFCsUDEtgpxA3CAm9+cAUN3j28n
se8ZShn1CCz9o8P2S2Gn6BzNjX0NYaCjd1ORZvxCksA36wvyc4al9bJvXFETKVv/lCQEbbqswiyY
PUqzuhdniWI3p5EwtJZVqsrYqNf1v+3rP6cholqfCD1x6Q8u2ZbSj1nite769YYbO+CE8OonRUTH
2BIOIi1pAG1d2Z+JFlJ3HnHKZttsfSk5QACtgn/ZLnz+o8gF150rb4gKOBco44Xfb7CRvgZBuDP2
8OOi6uNHEgBqo6jNCX+VycoO1LFptSSDf183lTF8/RS17HX9RHDKeuPUp6bwfg7ewKgAT7ZN0x4r
gkl5s5B42kxRBQUflfot4BshO1+FeVqO7NHXTL0JpU+JTxjgUMS/ViYcO1H7YvjFeJTynAdWLFks
SVWLLbq92M8RDANuoXgu7xg3B8qLuGQeWChL06Za/1cheasxiq8s/a8xahgGZG7DfIfhbN60HPFQ
McrbZPyfJgAH/3yrHVKzNUW0qUUhedVGZhPzhEslq/b4tSboOMxVO+DVsP+FW3dBF+07G/Yfc33Q
FD5P3blSxpC0hmBEbahAhDOTiLh4s0sK8oNN/7Gp/Xwdngv9tVltZ2ZjbKF2GVC9DsQlPjtuHu9k
/6oTRTKIRkMBrbY5qeHflI6cBsb7jYrmHxEUqkMwbt93C39m+9mW46iMCLEiTRHpnrLUS6ezDQOx
/LpuACgnU8BWz3/0Web4B++bUoDa+0q7Hcvr7WISnYPISSsOCFHAn74IWi2E3VkddSf7cry7xOBl
ijCI4ybVi2jTlFyYySR9eZpl1qoA6MVuub0AejD9PlKrCXBmPQpafSHOjzUdDzQg3tKpGtZeoXtb
LHPKBWd53xr82F8+qOI8Z7n2RhH4v4dgXbwTdHgk1DaGdEcf2wmdyiReCnXhQK+iVYcECFibuI35
ARe2jiteg+AimOXzkWw1Dy3G/nbJB5afqvIuOEf4e5xKFtffo9tc90IA5BlgcIm4GFGfZnMNplEo
6fWR+DdautH/DtAaEOPA9PJsG9Y7bkqjUVJZOSySFh+7d6BEty49b65OPifcaGhLJCpryhUEIdXg
huzdB1/9yEMgWYZDZZK8ndvO275bxBHRY1rbxLibhSbGv3aUXRlJkhuLi9PyQK1ZgEgpv5TTKPbA
ZMMTsNT4XgFfMurA6I7MUwMp6UMTRHaY7zhh4oX0Ckvs9jJ7nzx6ufmGfal1ALtqUU4n7LjTVOor
KSeK87M6ntkQVjVuvsXQutrREwqQmhLJEZ3zb7V0PGB6k9PGJgN2fb6VlhXo2eg3V0HOmoeRXUsH
+xN6V0N+7QE1yMzy2m1fgIcpI/OAQb9kC6dwIfAZQDlssO/6Hd/X0P8xxv4s5P/HkWABtc1AhRXr
4RxuWAGVzUyNpdoJRHoHQW26WURS2RLF5J2lzoIVF5DlxqZCBlEmJSQQNdru+TAjhDYBDT07Ej73
b7d9PxU5ceBMj1R6DrkWXPW/jAgkAIYmgBaus8SMEkzpV8EX48WmI8+jY3GOm3Q2v0uyxSTd2l6z
9RHncNnAFnRGgYFXBFwINlJmKfF+TSSRZ4imoBNGj6kHowXh7YgdzLCQJQVz9SmZezmPFCSs5k8E
ngXFWnmfdiYDWDbIjmoSJTymVCsxfHCsOiWzA0JZJ7daYe+rfWsULQQ76li6RqEa8u8fUYsz3s18
jv+sxiNuohhduJc/CSrnIffQKr+adYU3OkphhB8/5Iu4Cry8rdRyqAOPENNJLZBvJPVsYdeao8jw
B8dG93bCCrxongMFy07lnDOJLj4kx7t1a9E1Hy03UPN4eUFXIzPjbtlFueNI7Ln5DaUgQK91DKE6
NP0sOUuPcre7LuDDYoOiJDeqofWDvsG7WhXRiub/c1N5iYxV7gRT1gvscbd+dvF2/w6rc0i8NCIT
+pOy2bOZkxJWHRbXFywO/EPHg1i6c/OKQaiwvRY1lfftSn/AUFQ4odAODiE8h7uBMvZGl2unsWiA
MOQ4audLiPLWv/Njw4+I65xMz6KApRZQ1xihYvPqZDNy5WQK4c1fzoD3jBnCcfWhp+suV+LbgG9G
dhUoku5n/uzug7bHh9isI0LeBV1+uSnLwzpvRW7kgbsFFoCtsdpiPVdDbnRs0mhKjIH37RMAnSWg
1ajUsLhKDZ+0TJL5RjJU85WFYyc8yNOOOVbUauc+SRPUIwrffp1hJi9McLycOPMsgS0et3nrTrue
gP2miKve7i+uVvkBlMDIvWaG67CWPPZIgVIftR2ONtNYipzpIKh5T/qYHtQAqdxetfKYQHqM2q96
pNLg4PJFEpZOOq0X19XEqE2ecZDrg9iEd9OEB/irP9NzlPhUn3qk3GRaB1NOI3HsBgkxptWPtR3F
KOL7nrylIC2Ks7aY0+mlfPFAuI79JdkyD7KwMfqdOZ1RVyquU0lWwZILU+Z/sMcR+nj3epD3Txw9
ilWrrZByi06z9UMyA1kfrROfE2rVorphr/kdCOIfUc9SkZw1QRjjMavP/Fbp2bGrJL/AzucF4kQ5
WvBY3kZAZQq5ZHVIG/bafDGOtWjgyIBRgk4JtGcwacvMgIbrBrWXwpCoS9WM+PW2LdQSlt7njOyJ
H9orF+IdsqwUXs/PeBKTvdRhGLRD2tF49RIvLr/1SY+R8hzOlcfdx6Z9YxkwvjnONMIeSV82LKNz
xodXRgac+hiRWF4XZngtUfh7sciox5np1/5WnOgZ2UmpN8R/Qh9ZJSdH4LkfqLKMId7X6XDzT8TR
NdSKTm6fvs6aH+26VrkrWvSmKy0hE6QdFsmHGfzmNKDBsGKghsN3TEi404cZIM7xB+gvIzyKheVR
V41qpvaubqzw79+qzbyu+ljeGzotcSz2c5VZjcf65jWjYHusuTEWCH4MYTlqnU6P4TGceFPzU6nj
HzjDRfxpCGGTk8BJOq8yTk80M4Wr4N8WdZ02cp81WMHHwIOeO/NXnsGKtOYrQ/WhxBJlYDqFJOha
LiY5/wSnB+o0vEvKIueHyEEG7l4vrEnv4ieKMlkh2wu8TNs38tuRzEflsATwzKm+B8CzkDhmh9Hh
cuVeTzBoBOcK+rjPy5Izmtxa/raDe27m9AFb2TuiCDcKdm/K3xURx4KP1QmcqhS6aNecEfNrQmq1
Kps/Tj5I+VAuMWFfXo92qW2Us9tIYBImeY6cyu/M7ukGPT0+GG5LNqbXbdyImXau4m2/cbr+nvxS
c9yWxwo9ds6fYkHImbgcKra9Gtt1QSzsrj7ju1HN93OxnzBhFDr9Jg7P3u2Y1t2aDt6GP6B/hUPt
A9MfFHC8STexc+mparwu5qjOuXYP2j2Wqxh/8lgKibyj43LBmDKqLOajiUpcUqH42jP7Bu6fqNp1
7KZuXXaz1eQSHboM0mJn0O/Sg/WWzTYDMUl/G7M5qCaNOdY5bGCtTOAHxEnBjH7ep1bIGTuNWFdr
9Uwrqrsr7HrhdAQ0+XJL8JiEwQOntgl34eQLQJXqJYanMW7rQZETm/f8Wfgmxrpl3cnMC76POCNt
eIU28hqqGsQx+OUshlasc8G6Jim3qvHHCZFZHiPzuP6NJkT3D0rg8L9HQdGBhg21B0BtwRyGWbIf
fC4NoQFuglQpCBk9ZE4nehJg6OKf+BaLutB9S7dLB5/R+7Dwi01/CJt43eknpW7sIN6ENTua2bV/
2rYEuuEuLGxl+9N+8PpNNuHqAIFak6rnF7jPD9+/COI0PJwew3etjmBD4/+gSSe8sHm/0JcK2E40
il9nu9P4YkCMveqyYE4YX2vlmD+Ljt1nH3YlQ25ylfx7t/8dIZcfKL3Irb3Qw2nYVvhwj5pY64na
CSQbUk0ivKlIY9vkkPzbIFBdsLkx+px6xGxJOgW98PEwF78FOA8ljaRfpGpNAonV1y2tSI/kEuMJ
HC1k4rUxNcf6K32DN94VwjI8Qbo4x3g8wms3tSB5mAkYQeC5dLQ0B7WT/8LLXPxsipD5WmQuZeS6
ykouQJjzY81hZSneU1wVHOw0XSj1MYpqACRXxPrgg9ezc7GE8vDKvG35GDJfKJoo43uymQOflPsu
pnTwvqhDQjJrExRsD8wMIYk0jVP3X+KEoaVSyd9Hc1+nj+KuimAeqGRYNYI395kByrfdLgIxA66M
2A0KDMveTQ0EBSqEDMAPKsQHGYGwZ/gX/Y6Zw13lEiH2b8WkZab+rggW42oMnVr01ApO3cSKnMlV
ghhmNXVoTPRCH+3Qz97ZqLm/s0MC580JCQsrp5Ka5JLxMMsZ7f3dB4rA9khOgtzaKgBi7vEm6RCT
4haSyT8Wrp8hajg9yTlxKPzhUDJJr+SnQNx42wj+G7s6fpE7ulJykh4OOk6ABQ0vmGW6LdgBLSJV
DBFraUjGj18Izi8QKzN+QmbJU4ukC7tEBkuW2JuQrzAxprV8+nZIh4/11NrSmxLduMVOjRxS0bae
04rpqKvi2gN77Q09d695ddDAaaElCvrLfxKEn9JvpWQYGXrJd/e7eFETA3/ZOzZTZR7O1sQGjQiP
pzasOOHGjagRfh+ywp4ku791cWS1EZ7E9CXAml/qOYISYIDDLySmlgo96sq/XdVDnH5yr8d0nTC1
WcpdOY53CIiw7DJ0BojB3aZrXUswvzU2pPXaAF5E1819Jeao0UDGF8hzT91nuF1GcdV+GZY4Hlmr
zDyOde5PQ8S3XH8DbRVQMzb5UxwbkSBynhpqI6hiL+s+ws+eW2h5sk4BaMWv6ZmLoVJW8ujBLuoC
GFumSIdrK88jFqb0b5KLx83C5NAq4didz4mKA29G65XG9Yvf4+MKBFbsORf+pKjKmwodPkxeULqQ
gM+7kPXJpOcOFIWszxNV6CO5wKQngpuQz8O8CQqSieFw8QiaDNOc4J8IUaLOEunCHO1k+rhQFxYm
qb1lZThilR6jiFbrNiH4DsUz56BPE+AYiAMABjeAGpT1bSrzknv/Zw/sNrzsZ1oEnVVatpP2fJhQ
dnvtg2aJgRQi7YJCpH6PIDR8tMfYUyVm7Ez+x/1nndwi38kG/fn6MoXA991H/OBd8lBEyT8lKQ+4
Hu/cmetuOipfoaGXB00C61QeUiFjA+2y5IKOsWZiGM97Fz0sB2vvbDhiAcb/WMjWjRueMOHq2fiY
o48ndnTb4benUc2kOJAgObGpUz0O2UgSY0Ldnz7awbz84CKmta1q89MhK9AcWeCDQGQJyOWi+Fus
S/bUGeEKwltgDQsP2kGOeFK8GsW8NK0BFE2UN70jXw7N15Nefc2AexhYpiWd3+vv7tf0VbsmERPI
11suPiARUm24b61TuPsFiUa09QyQajzYO0ftlAlcKQyG//GLYOTu+XlJ5m6BHtw/uUYYWfVhGXT6
I9msygWspoc1vqR+VkgjGa4Cd3paWmWob6wjEQsWgbXCaMdF2MbPl9LFGup3VVG/CVWjyXZ29wtD
FIDIUuXOC+WzepPR3fB+o6aaWnYbvYC8WsFKUP11PAv0g3f4L0eZkb967Vj6em7VHfCIk6EomAu/
Exe6XOM1N2CqBbggk7uS+z9QN+m4J3fFEF2z4vkPRD+pXAoIAcMqg3EcF8dyzfHxO28+WUxFAGbd
VS3veyGmz49o5QwZsW51fiMPbbQ8ETtxpdZlsBu9z5cjFIAv8bNBazCN8ka4U4HLkl+zex1NBmjd
kCm55g+kmTEN34Hprt7/bIXPBpjDOuW8M1c+IdmY3Qf6LCJ7oudUJNf8kaWljHXtjevu772Zi+uK
tIYoaAn1IHrHkhJ19oaeQFMmmf1EyJCERvmWtKnGGeaXW8cbrZpfVKx4r88U1cACBzSzWDZIY3C7
PAzjs0A2CO9PT6Q4YXAIQnkXF7Knse0Lw1yIUYRuyQ+YZrlrh47imrTuYB6gpsrFeO0EC3bZZM6J
4YNkhS3A/mOX3LGurOR521b3O5EOJpGLMJTHnH/lYKtub29+Of8KQN2s8rcdkwUHTKwbRtbyszXk
rYzZcmjg5/rEGPdQD4wrqAAYb3YUjKg4umZNOFfEgBSf993Xry23+a43T/wqeqFTvinMzG/W6BcA
0w9Z/9vKDQLOTb+FJgFj6X7hKrWZcwkGTg3xbfuVqaL36TOutny1U9qXMepubcKxIOSM0TUjS6tS
D6OP1MIRl/rJs30NBKLseMlIlgogx5n0bYY5e2f/eA1lGbmjVXLLtKc0SCu1Hnjp2g3pMJH0ItES
oKSMxE7bZxvXF6pz4ivhZwn3sIxPA4uywXhWHDquWuZCp5293bXVI4+PiEa8HQoHqkZOqT8N5jXn
ZQWIBCbPbQ0Pl5Tp3l+Es/EIt82fpCAPV3X2scCrxgR2VYffRkTm1Vmnh8Fb/926q6Ds6h2ifV5V
c5CliLP8jYmbPuhOWkPZP8hgq/KDSzdFg8m7hjJLLwZffdk6SV5/8Z2o9mn6r6NduX2BC19c237w
5j+42wohcmG24haqpldZJma6vWre1T6SDIxQridWqUqTyuClcuFFmWRJ7/JYdwL/Fw0M4TYh4Zww
zrah8y5YYXLdOGDTSN6nfTvpoXox48gLDqpxXyb4NEo5V/mQDpDFghojEKB1OPtrT2/0z7uUXJYX
N4+JtGG/Xmd5nQFtxqtJSiVcIDJJhejl+iGpkchps7uv1RKU337qlPWBo0BlOCwhmMD3wqXkg5KN
LQBbQJYZKXRLzsoFH98iM1i2jeZYVnfLP4pQgKQPCfl3JEyGcSQaBl3hv+O4A7PtNT6EGzZBvJEg
IUcOwa/iKUKMvqLwed99Ml9URnEAkQT5KWMSiDe9wBn8yfxiuf2WTRlbTbFIQTS6VfY5ILJRcS08
A397QYr0pieuEE0F88NpDhWEF/QHRxBSWaO4aHX4X+hgvnB7noTlE2LvCINUz22MZA3+3m0ImxX9
tvz+grug4nxQn0HZ4pgTDu3/69tZuZAdgboOYly1/kHZTUKqENijF85ODcxqGC0s2Pqfb4yhRgS7
6wGT2AaP7pov6c8FCzOf+ulmkOZm5aBO7KWunKcACb5IDy7JcQOqzmI5y2ieFrutHCT9CMF5gL70
kwduFsfVnxQ+oHenqyP/XZDboptSD7HQQ8LRE4YBZAeQzvSrsG0sjOWmLKD8IGeCW8Kax0tgzDz0
55+cyiGT28DBO1sAUoojJnsXd7aBZmwGaUWDco1vRhkfURxyJSZ6KjWNHR48Do7P/OCfj7XRlUQG
WOnwi5d0dlvkMbumj+KN8Ft66AWok3Lq7FKE1gtLm3xJjhIwsSyu5jRDUuAioxeIaH1by7k8Qh3A
RCFEiTOdNh7BvGhmPPJLZraZIwGfCJE0nshM9GzMgr70xj0ydSGIAD8OWrowYP5ruKT3fjsOsmWE
wM6Knluhepmlm/i1frSLTzxjw1dHQ4X/OAtI2/3QZroPk3wULFkbk1dQvYkKC6X6tF9t4z1ywCej
28v9hPjeRYPebxeX/r8R2CcBgg/fLqSwxRUw6U+Go1yON45cqTKcw2CVWXkrVxA8vigjyDz/Ud83
SsZVKuNhnC+nLv16ykJN/GMZJNxYCfjDa5ku/Eh2qh/rWSRXb6T8Z3ZmQws7VSTPqQ22fiwbb3+v
keHktlnI7CkCEfGcYjNU1acJWVHrDm8d3RinUU9iWKkp7BUD/8Eirrg5kJR/GfdbTv1XZYBOozrN
PADVsWtNSF/4WKOD6xUacq3HGeiHsGhw+IP+p5m/vsRyV1MNMbgfyHvQe++n8Dv+ytgSmWlO6DG+
8b9dNBRedCJqWoz58xotnGh3X7ZsOzua6tKQODZQzM3mUG/ZnaOwrtdSyfMy2txXXOTyF2jkr0qh
UR1MLx1oqv6vjLLM+IZyf7OG9qBOfBtzkV3PQX+Z+nL9cWfZd+nOvgujib9DY0Kg7AdIc2xCUIgG
1WtLJgxb//gGC8ohfipOzIu1yzQyWY4hu8qro4wkF+3Nvb3pT6Fgl5JV/9Au1UVXzLMuN4trPoXz
f59BnpdYG7WpnPPv/MelvINp2U3uUdVyK9mc+mfpxI2V2qlBqqfEN/PnHhMCA52scuLoqnZ3TSYr
YR6BJeRPmVRuWnqx7efY3GlcfvUvmEHXFnrltfOGXTC85VXsGrv1KTjZcOTHo7QMhS82lOj7Z61O
c2sVG/wErjpBAR5+4wLUsfq/9JjDsF2gGxAjrbvHWhw1IeGH+YMErkdM3WrFE4CSDcrIx9oQzH1w
bRWtLTRu1zZFsQz6OUUBb1vqNBmcumAe/nd07URNxh52Py0mltHAvHM3epwTaX4K+UqHf5DR2rM4
T7XABmdvY1VRNWVbd6nI3Wwi+3OybaOE3rgIhUrrB/K9Pj35AM79v6CfS2cqlrPr3Ur0AukPlluX
EPRcSuu5kC2HBqW2Q1JbiNtFFzkR7frpxFfcdAprjQqgwglJhxJr5WI/a0PsGaPv1F4e6fXbVW61
GIVI9AdQULNTfMd5zmwNqxxFcIXgiO3416ZY1wtNajgSTdRe5mMzEvd0sCYg0cMbC+BY4lf77Ghp
y6yF/ih3rfhAiCD48rf6g0B1uT1W+1XjQkfuFAXUtxtBck55lZl2Wk++gIT12ZBgqRhxA3ZBvINY
WKERsAJMdTjy1N0RACJrsbNGdW/Eyab3BH+Z0a3vaMsblZgDQP4wM369KFY6LCmY6i5Qg/9TO1z2
+CIFFjVZi0BI+GhFKPJCToQno8WEqXXm3TZDcBcrwJ3mtZd4aQ2maHJEGSEn6cf+/QUeYJsgQyDU
39pib2CpctdHfNWb7/MbXDR401MTCUggimjej7pHywZ249ByLGxQfWBDKY82vMUyF9Pgvx4QdlAa
arWbgJ72OJaQ0d3SneBG9Yq8Es8W+yRiLQ3t2YSJsRB1omjUEGbZCUSqsW8a6HjwnqlZqLuhMtyx
G+XjftkvLpWWTNEZwIfAT8YgsQgdNsGn7Xk6OD6N9W8CFCmrLaeNTYgZEYH99JLxAXNIQHCd0zHJ
CSmIOCLB96c3gOBwM8yB5zWv7E9ibk5sYvjYADL/ga3NPlVhoAPzzSx+hwfcmaBgBcSavO6DfaSz
ObXEsgR4rkfwRuvcJb1caTnJEPYcObVGIZEOG8MettI6EmZ9Ap05iLt3Qla1/n0EXmKuiYe+wgum
NVszR52EdCyfNbB1gj0a8wKf8u/4lM6sQ1xCthVDNZnHG7IbI/Yqro5GgdDRN+gUbYRZFp+8UmHB
W3q1c36N9fnYUvveXoLCdOB7KMEMdlqXKpIUwQIk3RJFLr+UXOnmR8pfPRf34f/KcafcIXFELeC+
zr6qZoaQeSHYheY0Tzphe6lbEVN4zH4Vpc2qxuij4BokYOoZnzqatAv1KiCQIIQll7GeEG/ZJVCU
lVJ5qxmfCiR2k95BGDbsI70hwxXs4A4HKVjUtiCVQpqrYC3Drj1bZyBEEm/Zuu245WLUaoNfJ5ib
8RPRN2UBDnxlNc5GjH4wBc5C5cVO4NhsDZqAJTn2ua1lbydF6FiyVVf3aufwK9LVC287Hu0JrolD
roVA6gmVpVzXYJMxgq5v/6V/e94VUQNwcsFmNeU5YroRONSZPbwwWA0eqnpYNyfsKnsNNi5QpOVc
vVhGD5wcGNqo9S/pFCZL2bpHnQcB2+RNPIdh/AuybMgulXc5VbflFTSn5qblHWlcikBR7soXxaIU
VZoDE5i+SzatvwceBy3zuxwHy2T0f8VBdWx2siOWLDUJgeRfW9z7W43QozecCL3BrTKFz4rVkbf3
vwPQ7kEI4fx7xrsKjbeNfgFk6lFdXWn7n8JIIb6DZIFvD4g1EYCuOqNUd0kvI6mYBKHAPRYsHMvY
XxIwQR0juN15RC/TRUXPpyphMSleMdNOdqVPRCldq7VrnHS0ztC22SQ9wdya4EURLsJ1h7NM+wnw
sX0Ansps8vxgn9Y8R0Y7vx9XaQa55VM3mpKd9835J9fMZGazhL6VGY9sJsWuLN+SZc1K4x6qIQON
IaO+6sKQ4V7GKahFbYHRd8HDb63Kyyw/KMvyMElIe3W2SOzhwS5jemY7iyBaPewJssmJ8L+1lLrE
FPnApB0Ck4GcCinxCnseMThvY+/WHpnQvj5a/v3hfPYTsRArb0fqgBBZtw4WL2KwjW6DF+X3EsAn
3fj6nocC3dDicd0qQLld+KhZP5jWlX/CToc4RcAEIc+HT+LM7PS4IyXUiQQLd9DDWCUrANAVoM0p
Z/2kdpEvEIQu5XUzmG9CfMr/WqNkOBN5lu8bm/LqnaL5bAk1bGNq+C+tf1UsR6im1yoZs6kiCb8l
nZLD2p9ZA926GJUAsRiRH5ySZwpafhcpfCBcRCE9YilR8fIzw/F9EwEbmHCgbpZycoiO28L5sx+f
DDX1iR0GvvAuGLe4lfthxj+7GKkfCx8cmBlJnYfIeMj0mOh1b1kUU2zZf0NwSwVlBqAMXAyh1hol
GBX2m23ZnRsIVv65hvdPhT+1GWZbeTs+pU+P9/Tsm0OAYnbNccyfePNFihzuqueQUGqrYyURWYzG
OiRlpATvFskSOhW8zgwb5uhmGQAwi+6jIh514wOhYinoh7WaSGgrv5n/PUfJuzZkOWQtJuIJGBks
n7Ht7vXNVyl81yZ9uAD3/VNyC/N0lZLDjTTp/0VXub9mcfzJFNWSbKXZek/MtBQOS7weHNNhwRq+
lrBDepz6TECg98abAg8yOamwdPDRLEKzlQtVNFRqWcNmJAn+O5Fkt6EYvrS2Mekz17uIRomLC/uh
aKNILavXO43fijr2siGX1LHipYTvjy917y5vGGKhMvERUrssFUrksukeA2grbcJvybiCnTAIXYqZ
k/5lvQHO9QSIk1h6h/pJi+SCEFCRg6RbrEro9VOoTk9hFEgHjReuSq8Ax3xf3ulXWTvnCeRJH0MO
DOicClY4qVmrNpQ5Cc/hl71QhZmwBJC5VRsEEUqG4J6P2FBIDVDe1zNORedZcLuAZ4UQXdmiDJcR
cemfLGXa3AeaeKBTZ60Dp0qLHVxK2hZgz+TPEPPFT6xq5Ns29PvZ9FBQmL9qkQ2fut6J9lwqrssD
eSJrkXoZ1oIfoFf4+PKXaC5jQ/4Rfwfut9wQgpJ1Bc5j7OqrRNQeXig4veAH/4IsPIV2x2VYeXV/
2eH5f8VAD4hLajB+yatPK1h4KWb6Tbphbov642JqQFhFYH/9bqZ7OPE3NROtf3ceg5ffnFFoyFpo
zSRlt6vn+aZS3CHQojw9U1X0GsHP533naHZmcTHHLafyEbjXELHNNuisUZ0PXZOQpUYh/gcU4r4w
W9cIIHoPgFDG8GYUN3EECXCbzgPvBNZIOYc8ey+6yH5rbBE5j4bBMrWAD/1eSMc77EGnrWuAViqp
uFY7WKp2YxrCa28qgIqhycuqA7/V44WSt/c4KLWW4N2yz3brm2KD0J8fyiC6FDdfk8cQic+TcdB7
ntNlxXjZ+tCtvasHC+SGK659Fp+9Jx9K0s55Uu3ip+hAIVT/72Kbxyf/vDIDSJeCnXbD8co5RNq7
4AHaDEfq4nGsnTWJZzTB9HXmZWirsfmUFt7fYrZfllVQQxookWWCfORy6qDhOf6t1WU7JEWqzqt8
HCOUL5+G8+W/MIZQHUKeGYhXCHPsyDzFkwXcm0lJ++bt2mxmFCudEtZ9r5TYQzcuuDkPC8O7/r1u
JjHz67JM34jkWCx8GDAmS4OMmcA5id9EX27J/S8cpSF4OtM1vZf8dkb3iAV9SMIF5iJ9rNzpDe4l
WqE7npRs5BzJ0X/NFTR8VPvdoIQDC3RjtuLcd3Pa5VZxOD1vjpFrV8EwWBbLflpzNGjhuNEv7jbG
ugahqRNe6oQluxRIcaaM3DY6KbPyi7gmo8B5cw6C1szDZR9XUvEC5ciTsjpIH3+U+BMHOB5l4k2V
qFzilMYS25WteyU1D0MrDxX5WNbmM2oJCTzoqD/HtEKS9EqkY98kxfH7FZWI5GNzke+1qzfXf/HE
kMlYlP/N1DVwTUekiPiPNwh/GldnubtGKNun0+i6eRivJt5fYXvPIHP7kvJnbsOUQ7Lwbi/LWvcX
fEmn/MqMlHH0DM/1H1h3uZCLgeIC/ecUv5cnyOYPnx4OAajpJiD3zUlVBuhDz48UdCth6y0q4V8q
c1RYF23C0+xro1RMBi+iUlhoQbN1uM5AMTRSFtpaRR44IxebICQU/MD21fGoOvO1zNVtmTSn1Mhv
oY7hR7rPvZGvVy7ddtzqR93Fsf57ww1Df4vS2kTuKa8eideEOA+ZqzhAOxOuBKbI0vRfeaNoLEk1
R53+RtgoreOOWhAF+xz/1FDI59RoDFs0hZLGYsa4bVz+LtiN2y/Vs+hWd+Ab/Cwm9vBpoJeGxHZT
QmEk8dF77RY/8fuk4KS+mERM6q94C4BK/+NB1YZtqcLMhbCsNzjNaJAbmsOCD5eBaB1BiviP6nwU
lZVvyI74OnfvCRfd73Skwn8/BKTiLjB+9ca7zulwU0iNdH7i55vzbb1/vQm3YWJ9Qfwu7g6FNtwZ
2aVI6UoCsWAD36YDjmjtiyQejs681C+e5+VneYc1YAcmILXmjPWwl6j0wZMLjFE+7SEO5OLTz77J
MrpGl/SeVwXfTpbuuPcwrMH5OzQIl93CmsHmgw1Z0OMLITV1pmLEL3kyhCTSh4PYIWp/KW+JhNw6
vPRVJY8P4uFKfhfWvI2pQ+3ksY09Z8POvceBKLGusGyq1A0c9XwVmC+xLUxsg1qU1UHvkxnzDU+c
aNParVbBVsso02O01Az/hbMHfEFjz3yex1zKky8ZPj9wtuVSwiXZrgF5lpmSoTaMirJCuKC4tc1C
J2AVodmrqFG6ZvtcuppUIi0qZywmXb9fpif3/Quselvq8qb4r2RtuhSe1RT5S/+gGAar+6NEQoiU
5aqNIzTOIaSvNnvSN/xl8FZ468rZX3gyDuqmWyg1DjFc1wGBopA+Mo8RhSzru2X5eMZXDpWPsx0/
xKu/ZI0dRwQXxK43iof8Tmg+2qzyTMjk4YH6FD+lXdQgpyWrGJJFVumfE9GU+9EdlNp9EO8dKJzT
XrTY9LmtYwR2Mwp1pG+E0U/nwf8xjC7xJwKgYR6GwW2D8OK3koYKClC7D+U70vZiUh+POj4c8b73
fQrT+rHPriAR1ybpcKjgrV0wdMdxPGZkWbBByTpAOgli93iFHPB77qVi2idEfEAjwPeZhSeG2KDC
ShX+5Ljohi5VPifAdyluqPAIzL/qxVxOSF6qkMt5p/+RCoh/XW1iJmPrAdESDJt3fYuQSHxS/qkd
xbhhqN7GUU3Wg3OrudbgRCiMbbIY0Y8H4/eQIGZ0/R7aE2YGZ5PFidW8z9HoqXoqPPjQDQHD+w5C
tPpZDWxD4SAL6gOWw6sb2EEjt33+kQjCDbd1bYn90I/8cyXL1GktGaNHaCS0VpRWEw4YxaMLFsvt
BBy8dGGG/TQB/T667p5bJzjWLSUaAgpDiVxmsD5hquCpQaYxpVbrRfvE3XgAmUnmlTJqZSQxm/kf
Gc6bm370FaQpwTjFLyYSm8TgQLI9vXmS8GNXqmgHRsD1clFv5i4fR9/t5vBA1sJ9/7P9dSW3Eb+H
jicR/7gbHJ9aFWBeAX2MIboCgmEqRezQajzW07pdylp4a1rC6Wrw+ceGg5Ndkp5h4eY6RvzvePUg
EXcTtai2fO47Zof6Rccovrwhb3yneDq0XqALF0yS+IXR7orrwpoU9R1yinzkeO4gXIYfJEGJUUm9
yjFtatQ2R4FP8wqNwwosi8+anspo/D4FeqwxioxpEglUsSiSsSi23i46dFfRJ9DOk/dh7BOmh1vh
ajUYrpZ/Q5d38WX8regp4rhk40XXcXP71eP43zbE6hXrLBaHQniQSZCyB5lU0cHMhzBxyXcYSGHc
++4lAdpdN5RSrHj1MSXsnN9X/zucjxqNYZnQEMADpKm//G13ULgqXIyLzc4V99b/6T/iFAWyaNne
PCi7x3dUqMogB73PtPnqGYKQ++zQiLtQhhzRY2Jjn1+RZQvgcM07FOW4K80KGYLM4AXL2brDHpCL
pR/V1TeDXRUfR/OUEVBwgUr1eh9Zjao3Mz+DzKEn8Z1IUoyW+MLRQkKmOFNxocG8RSv/aynJnD8D
mVxWkvX/00GpA7ldYp6LeApusODuPvc5zHBwchWNHyK6ma3Q0TR05n10cvsAljczzVck266CYBAt
k9aT5fX+itGT+/Yc0WMW9huj4GiMy+EzytTeSLjamVmU9wbUB1vPO7ct9BrahIIAl2gogvhOr0nB
17aoqoPw4rcQPontYBWLpdEifsUFLCwSDMZVmn5iTdSgM32cPgVThenFJ0+cSp6reH8BbPnkq1Hs
YcXfURZ4Jw59Juuz9ie/STvAV22UKSHkXTOZIhiTzninK+h2UM+6vGEstmC3R+FF8VU0SoCprIuw
StXsDz/z4cJv72EOD7Ru+fW5upxtTxFPmDZcexWPwUADWLp/EECr4cWf+kSms+f+pUhnM+zVmWES
oLU94c0OSjZ4GkRwHJ0RAQnWN2sTVXTi2xhwUnEdT7TaAmMkzDEwfrI48jT8LZ8sYfjNpP7fOeIU
AEML3obpP7GO+dCXfR5+Cm2rRdb42ytevboLA/mXpSttouCxTUkPOCVkR8dbq2rJkUjYQ/nPz1p5
MsiPIgW+P2yCcM0F35YTMwKnn9g/5OOQunNoorytzp/Ez22ojfqCfe+gXkclTlxPQMEWRYIjUu4E
Etdb6fxj449o0CTA+95HqkSwPsIKr5S743EPL/FfTEoHOYA44Y4ySfeeqzSzqZVGzzEjwBIS/tKC
+QWNSB+mCMx9RtHnhvmghOdTRU2KEsjg4EzlGXWUodnrTu7vIT79WQmotwEpXWBpGeSL9YubfOgh
Aiv6DXQ31hAVc+5Nq0zWOMdyU9tGG8PoI4sG9UiDOoOd1JokWLKSoBuFef3EYg+8cuWDHp/8aUhh
pLTK8Zi6hhTkaZdPLRRDLrZQWCI0mfo+77U9H66j42cmtSUP5estodc1TOegintCdI03/tGAaYpG
zKs35w641zV312YdtDkAc138SVMqL+Hyjlzmk4qThffJuJu3W2uuVoWXTBBe/fKo8JAQ0jTNsndx
I6Du4p7BYyU6MBiBVVNf5+Dx9BiH5KH3Gey5Mcd6DaMzQHv/A1hbVA+IIF95axAdq6MxP4SQOeH5
7VZTdwGi4R06lcXNrgkPqsK2kvHqf98c2/FJpdJ0CjW0s8V/AKgi67cb4SG5f8wdfWLSRr6nhYpl
RmvEH3QoaOBkArUnjFnnoTptyWhMPLootLxU0bzFdnNNF5il+gK5FMPv4pCo5dmIqsnJ7T5Vr04Y
ELzQvQ9XmpXNcbFZAEnSmZScVIHCzJhsq0yynFYr2PTz2lzLjTEXvQXzFjXLlXiV+Yg7GDlLKxDx
12oboD5nB+ckz877kMaX/n6WpuNQWDfI/8E0KTWNU+TgAD0ycXE+m6GvMiZQD1JWcI2nqvpJeDSp
Io4H7f58aKLUG0q3MdaROoT1O5GBc0Aqk/kmNuHQY4s1sxZ/7bbVqV8v+VtA2xZlIKfqxaz8e0uG
AQ+5GBgZVArTUSFxa5+gQxjCyj8pP/8EobkC3uLgy5kg9qecU4grOGoQzgURbk+mHH02HOf1AhA6
o63iWiY9jzuYFzx3icxJ9d6UlXx0fGBu4cwXKw+fo3+kHg6DJ01kP/lrNdh6meza+hCBKGNytaxL
jBIDuiISjOAus3yc1xrgzF5Le8zVFWh9z8Lk3Ce+1A1Cqnb2EgHXAo6ho3rruiFkTs6wqi/xadFg
WhPt7mmGMnkBHZFeIsKwYEzdzOgTACEPvcJOueO6FrC4o5w61NKh2PjlR+wDIXps39QCrZw92dHi
V9aYm9ePZTcLnEMbqW/Obtxwjm+WvzjqLOwKZjNljA0hzDIJV9zCqRV/55PtI5/zV2nqW4+DboOZ
1mLT2nWj4qAjaL/iVNmG69nGsojaxDD/ht0vHrMI6Bs16wlYx565DYa+QbBSw8tfjj5H6dyKmpXS
9CZXvzJRrJTahqJLEkYQQuju8OGPOLIY8EqRpnGe+hheTeq00phQ+0Zz37O+5tq/3jmZU4djCe4o
g/ogKfd/bXs1VzMPLE5Xarh8I85JSlOduVHFPOtuREd5ZIi2+zdg2XgYgYwX5K80CyH4byhEKwaW
3i8Qm3uKmAicg2CW6mPTPJy15fFNrH35TIs2AHWoWsPGOzeS/Eb/J1vrVuG6kkhRZkv8+2VF+TXa
hK8Mk1mPuOXjrdmgZMkZvzTGOHMVbkH4DVATgnlgrqGG7TiKzFUdow3jaAXhjRwg7WaNECQmQva3
AU1D80Kf6+BDZ8faPQ+l2AC91MeUceKMiJ4/sWgyvfzPdmHGK+AlyEF6v2yaJ6iLBcusVwvzDZOR
B+1JjNUwYfxpC+oYPfQXG8KC9rSEaA624LIfOX1N2ZNwpTMcSczr/poQzrB9Aqh3Ymg5fbgbFHgO
MMmyPDgM+qRU0JIrMjnanWVorjJuTLB54fmgTJgSJEgf71Y4VgWPO+NtQjUL9gYcMzaLc5xE1Jiw
sJAEkxTAUUDcHk4d0qi8iWSEUSRFvDTUpA4V3s+4z+LYH64ud/5lPYMSNakiOC3SSaNanNdDnrsw
TXG9hMiLuhGa5NXtwKJd7G1smgDAWKcWrYO6V1+KfZRehAsYcvu/fo5v7vOHs8GliXygESOm7vk5
BiuWq0sJmQkiTx8xf/1oN4g4GlzDod2DsiyrbM8T8PO2YjnrZOz8/lbd7n/3Kq1YR2WWG03dfL3j
frycgVcufZOWhSOJD7HEhgCd9dJhuLRQTzeadUMfwUqgOfi/aCIK/A5ZzRy9QF7hUd4xzC59KMc3
iNRufuvwGnCFFLDArCM9R7HwD93XVf8xiZZ3gglXCStwgSkYM8SBZZ/kj5AFjb8DK0aNVIOOUYAk
X6RDVccGWEymBKL4Nc0iWYeojhdesiqjic9KA9VM/X4lOW32ZnSuCTgnVJIN03VduJfeIbN/QGW0
1Iv1mCqOO6BHIoLdI+HqhDhXDdPOUGwDcIUGsVsaqPC3jdxjZVpWsGHzSVTdrA0TVBzBS5nwfjp9
OYe4wg5g1bm/BaLXAXJJsA7WUzhY7JjocBAuzAw4IvjEdRVeAECwqtNZffOsXL+WzPsNFfT2p/cU
PedluF8knHeL74XCtvdVqCr7D1aZn6GQ5Lf6JmxRybd2OV7/Zwh84j24lqU326vrXTzyqEEM48x6
NgJLmWqCWn8tTgl7+WEKk/UIHRF7obtsPGDE/OzDAPILN50t8+0gJdo8VONGT4Ew3N4vSbdSVnaV
kUk1MCjCwlzmR4Vwvy1SfD3xLknu3PgdQy1/1EibUhaKzlhfIf5DsZ6RTMiHWtuYKu2782dnzPGM
qSMHfhITztLG8pg07ruH299Xj6uRS7oO2H+/alst0VVN3La/L3yeVrmkg+KeE4mDodNEpeciHkp9
xEoaWaMXToFUFc7m1pN9evWG0XcVk6x2PlLrkxpThPfLVhS39wkI+bUomkebUxA7YwO9MDrrThZ5
741/IZW5hqifYFc3LYXcaeuI47C8GXNyW57pGKl0oUUlcz3P9XGhXB2226V4O2reobEUntgiXJhQ
KsL30RxxLJQONsn1A6H2csOouhrZYInGLovs7zQz/Nm+YX+EJ4ukqV3wrxRmKAq2CYvtfzs5nYnI
1Lr1bHMIqexJeRissnCALoF8awpd/D6/QcKlx1zqqoShVfPC/ZtGLIEnAATNLVbsorpCcX/ZXz+q
BbZyJTUVnRm++Jyb5maSUxp0ksxWRF5R6RJdnWcx3CzWYfPAD/wvXAlv5waorrflE2MgT5kRA1IQ
jHe3o4JHcXQd33TR+2bYo8Jkwtv5tKyEMdwFKtKhlpA11CUhNzD2zFkQ+iyIKmZinEAsCSlvwKpq
ma6wdiHkVB3KCmRFm3GUU8FQbIHgRGH1S5LVJKy1Z32UHZ2NZEVCn0mZk+hJQHGVfYtuwtAv8uhD
zkI+XHgRC94UPWtPxq37vdE6kN1L7SDVap45n3rFMaJRtkbu1aMr4OC4AYeN7O6eh/WlksfE9EAJ
mpPI3qhJFrvJuXaxf5wCngPqOkEgIot1jC+3BorV0H85EgejbY6lSpBjtVResnBl0b7l9Zx43/HO
W94I+GM4pdFktedCSJ8+X8y3aEJNBiqPN8aMG6azxI50DsOg7vgX+wk73Drlv+Tl/DieHA0bOzCq
oCMgYCv2mxoKv5zXO6MACya/EeMu6jR6VMzV9JcXEjRk19iP/BePt0VV3INRGut97dA83VEXHYwo
qNB5qcRUhXJokdUnSba3R4wycuo/GssulNqkIZmP8ZmNvqjv2VTSHCEr51VbNeeZwXj5QCEfvkeh
5IO16cqR82tZq8RKhMkFqgllVWt7Pl3fc6UJGMp73znjWu9BwymZ+34YiyIfvO/eTZVb1ClwkYCp
/+sNro64iB0dObRD3Ceud3FEdvJNajmjfH8TWnVLp6AF2inRAU8EXT3WsdLqjvhm6EPTH6uZUMUB
90KZvR7qVMINKE054yH+NQATx4CVpj7DbQLAjzaSbTa29TtBhvSTgMd+kMfrLDr+E4uxQ5J7exYX
+u4lZfrah6Q1L3PvGBZl99GBFayUKJpAYWwzbk7mjJnl445JpkASXhooe3V7CKyPQHH2u2S74HwE
z2Ron046ctGYnlK95gAGMM06XSC42fXJxfh8ss6DVHtaGf+EA6AzzugQmRRH4GmDpr0f7yUywTzt
ldmVCb7DX7vCDPtkPwL8+S6npDklfO0Brgi9C9dwxiRus5F1obTUbwT5B8swp5BMyEm0B6QoR3TN
a45wu8vmRvKX/+rYzQ9Uh7cv0I0qPsbh/CEEvDFHPisRHP1HlQ2XYue8NItjJUba8mmloUUcqhEU
QomX+c21ZU/cRhUkEZ9L8XHazixAn7aNbgQGb17uNJbZjsMrvrxR0xwbEdeAIQPYIFQ8HSY7feKR
80LJY/49CRgL4VAcx9NQqM1x+o4cjkunDCAfQF304SbSuWewCeVVqEJi9obzNIWtKXM4ycFqBXdJ
0Iwa87Ql2zGXt8ySxEgNOjmbEh/u5EL6NXOp9GV5hmPmWQBk2+w1hnsEGwOoRv3svt5DtoQYIO+z
VPhlYPzXROjyFQ+JNcWWddsIGMf8ueIhy0UvkNALKq56QM2IgHUTQ6grWcU6lJ7GdWJvZCvbL2tW
14Thv6qmWwEXjmXo2XnI8LLY9XHhYb2ws6ql6Wyn0kVnMoP27ctEhymYRGSIeYHAwIDj+MlfWM/B
TLhuxjc1i2SuSum7Bn+LCTThmIvXcqgZEDwD8KtBpsLN+Jd4I7GeFCDajLX/vEffqk5KgnbQL21W
XCQtpvCEZUTC1XnUEJjwIJ7CMuwYXCgMNyhHWRgH93L5wrt4P1e4cG9Zn6184wVN2dF4VmP+8QrC
8yX4OvS5ARQmv1D7xqExkHIyeAUXx9ES9vmB+5qkxfSWTIvNioLwp5KVNHvRb8R0mePwqK4zkbJB
bqLOTvDKDHwCqi40J3+s6PMxzKG7IKeyywhuBRbaqUwIX9JeFr29RgTelBovz2Msya/zFR7Uq/nO
hdsWxwJH/Kxih2tBFGENc8yf6apgbGgJPc6PRWShjqZE4Om84ZEDuDoAAPXM6qPNcEj9hopqy7rW
S5N9cBgrFhmFVMmGQ1bXANKY9g+G5obTKwkObz34Z5nem1HKaI+3WGTNuxd8/z7TtL2LQiV+sIy9
9D7qT9ryq1xgKfhWeHRAv9Z4ostGkD4eyg6SMVuy+W1rP/dpH77ALtR3cIgyszh3e+Iumb2J2iX1
nm1DvFbcZVHr9+ZsrWGg9Riwu0Y4JqtoMioUIOFElSBVQWkl/cFU44AsI8MkXkhPJXWp3lUjaSD+
0SmshFXmsNeRihOr6NlItLJ0DQPeTee4h01HE3G+Nq0nNXTLKNFOsZ96bVXPV+hy0jUwxFjLQzT9
BsopEEjiJnhU2bSq5o/qn+MugzmTa567oz4SOGPCGL7RmqKNZdtjJeTYizWdZNCbXGG8CVu3ACFB
JDYlKiHsob31pcfhg5qS5AMcCQcf0+fp2OCad6xoIYPgC0vFJo3GvVQv07uOF1MpC6h9dUt5hY3L
hQP0r6PqhLzaxmsiEzLgPvb+/V4bxDUM4DOQM8MTb8vFUyWg+YUPjhkrgt0wOJOryZWD4cIbWU21
TwCOQSfhwZgiN2WXbynUyRix02yh6fzzQJPjeVgrJik2Vfd4aQ/qvyEtyDsvCibsdK6/d59aRxcv
0S9m+8rK7LHlLKrLopFLcE07o+TxpZoAG18Si7ug9NCHW1Ld5yz4HwJaJBQh37Bhe5wmHDBDIHBF
9KjzWW3gHPm4LZqNyAix6yrfplcWtcLLB2Itv9amNzeyoiFTp6gLsy45q9K+TyDQya8rkTJqQFxu
xMpRYf4pOi/OkOeFD24ZMo6FoX2J+toc0bnnox8ZUTgC5qqEnrW7/P07/Yoe36/4fV10/K64sWfw
RYMb0wqPCgdemYyNEkqN/4TTCiMvFQv1nsKL57mX5hNWkZQayGQDhKAf0RWKC3I2CVnLVSysf/m9
9gVbED7XQDKzJXndiV82UtgqPOPsicP4mUK+WGQAOsHO1EUDNTPBehjIVEvCLyYKJYjwKiqDQjVq
iE8s8sKzVr4BkxWiXUfvp6ZJTRblFmWv202nzT3+NAxBp7Qcmr1ayf7Mbi+GK3U18qbsi2dGOXlK
1HCm6+jHiEnLbd/Tr9ElrxZTofzErkCVigU3NHdVAz0PrXyTCg77G8aBPwuKQTcFvvjTmmitiKzI
rCp6MTbnUHWl7QYN1B/yCNMnVLIdiWDifU0LBQDZdIZn2zC60TrPimnlZ8dkNk/9U/CSUZH3vDhZ
VtFPq/oClZhjoS8ISfIEsYyIMyyouCgJBfd1OfbS3uZW6hBWtqHBrST6cp8MI/OLoal7dqjNEnIV
YU1YDHgLfc0ohp5NNNOrkPF2HLL4iRDh9KgtoLRVSvbfkQ4TnGeCY2dvwBZNNBQYK67rGRfpVCLh
iyMKihAVCEMtXwf7LtF4kN86nVVOgBYiPdzV0wvvhHL30Fd6aDESe5o3mOqdT3gcub0+DMM4m94j
geCHhUxooDlvvtvPZg2FthTm2WBoejdSQGJQxPNuDcp2guouCqVPsTqOhMCkFa7B8VopV0ogsN5U
Iv17fCde1ILVOWqMtZcSo5uU/7R+8rAoWRmL5W2lY2xuHSSslCqtIUOJHRba5IiUBdAr2ffGcC6m
egakw7jOkUru3WO3lPToxAACpawcZdZOvGhZUs4W1GZxztQoIhuTDvmPJqZ0bEB2Q6TzO//0hEJB
Nry+4NwGSIq5s8bGRcUllkkCkyFsjSnbpTTaE4P4Zm5VpoAZ/Oe86vxs4t8898rMxtnSzMysvdbY
c19hgVsdMckuGaR7LE1DNDvAWWyswhYmTHJvGfqpf7YciWDX9Bbxzlmu5KFH19o6BHF+9iCSYkSW
WX4ZigrfgH/3sa79xdFfApW0TYkZ0Sw2vr+1cFlKqBpiBYbwujw1A7OsJ0tkoJIw3YM1hso0LXP9
L8pYvxoqdIoncmMudOXFafSTUlVD8RtOoKZ0bMfeuA6y77O+AThQPX3cnDAPNyLzonZACjWPuvFR
titSXctGCsr3vrEQBi0uKWe3O8GivKx0PIixdb00C+BQTfhjr2NNkv/cAyu5bj3Rb69K7By1e5ow
rPNU+9m0efZZUagC0+vgl00xeS5vno9NDcJMsMjq4CMf3kVpcZRLlUapBzlkbrJxXu/ZHuAJS5y/
u1lRmjhEY3kqzkUIvmpNREzi+B7/2TdKV3f9CwyUF3LitVtnAfMAunESSEh34Byfy4M99uI1Ai5l
DFxD9zvTyHwbuAvEy7hnZRLnQbWSLd0qVviXjUdoyd1Q8AwRvOPnKaxmn4Ti7Wrj3p8550asKcBc
GoKULjeddvD+sVLCejPt/qDiVysDM5UPxq75XAtIWUQU1tTHybXlQ3wtTss8+Y/O8LuZmjvL08kj
IqFB1c0a6tw68A1O3Ap5fnJ8enAgsZfykoAyn/LSHNu292kaJWaVXxHlGYRt1YKz7mC2XicVkD7K
TcfO39WNHChyi98QsWhv0YszWWndcolwPGk7BdJfeI7H3xWyXmZ0VIKAdkbR2El3mSF9C7SacGuh
BMljUba5Nx1DORYP9pvtUzyGn27TbQnpLMxRWulPuxeWL4Y1bXMNS4wyhJhCRO/IWkTHIhh8J5fX
LhwPQwvBKBx044j4SkGCYwvT6kr0vZj9G5Zx7DBJ1ELPJLkgQIt6t4NgYRy457IYIs9NLwvxxHJ1
MtTXyRZi9Ug6LWmqBpR6crvhUQbsoJqccYxXf5nfd8XMYNLJnVvCTY/ORNhiYAhXF1TYYL+iqSvp
gqpRBYX5XryOlDXkqfbREIjiebaEuOI08+gTy5HYXig2AMfkt0FeFh/nJHAFH689zb2yj57N+T7X
1UZTNZKaIerZcHg19qFV8Lnag0BlpGXV9YWQTuclCzm5m2sT2t5LX7c2x/7I7QH0eEitwoR1W6nA
SInEsUkronpdjT7QlEBsvqFJJidB1jM2xTLLeYqtRVacP/OW5SvOIoX2J7lLg0dEBtY9w2OgLnRm
sUDyEFhiJG8fMQQYtZq7gXduMbWJjs6yZxjQETbl/y1Li5gpRdtVMe5O+tsYl47tcBt8s7f5BdGL
gDsAYul1jCkg0Tp8x07falhjHkK34pe1Et/Ri1ojMQ8o+1w/moPwsf9b2+7pzu+pDaGgRhTFWYNJ
wKo1BTrjOHcu7BRCI23dnFHw0ecfyW/lzol4+VyuLIopFKmFg5OnlAkCEYpgBMkNBuEJUmrnlb0j
uSS9w18pmRI1XxufZQ+8Pd8VvIFD7+9WMlpP6QA90seUSjV2uNNKr84L48PVHbhGLOjQP6ndaQwt
cq7vriNkyP53hIKqP5YteABXGQxzBgSSzOnIHszg6D4HnDumDWL4fLvIiPcqB6GbtBImzZhtznJN
GwrKS+88+VZRJDEkHUKnHw9kB4tamd6I/C/IfUDTECcgvGYHBsIjWuI+AG4U8HGHA+Q7HVNy5i9F
0DdK2TObNuL7jwfEan1AJSCB2edP35P09V0iiXNWby/jrhRz4QY2P+JJanYBr7dHmMpml5fV3F+e
Gy2apyWNUYqH86sRVV8puayQbPyWDhjngr78sgdegcRGnlzsizDInvx49DcUKFECqEp1fq+fAe+w
mn1LXKChoDAD0kJ32ociXYtPxYpNQV3JdKgsIb/XSLamDnzfLfQa093Ar6+53OECrFsuWAK8erDw
cC/lKvrJ6Kp9JO3vrAmAwZXFGwPLYiOvS09BK8vPf8+c+cVkvQJrsNrxL4c7PskP5aCSIynjjlur
lYPdhqBpRuCym6J88SpQT4n9H3iwGBQ/zcYLT+lMSgsm2Vn+cPrI/YBAJ2b/qHR6yLGkUw6dQDgf
uzb6egVXbfmcTAqjlIwqnjkVB3wpBeiUjR04PFdugeaMfP9TsU5qLsLY+Mv7Gfhg1NXwhzWGmCOm
9UCZENpJyLURUJwt6DPnGgeYoN7ex30q7k+unnGj+kCvCrFqE48oiNUHG5FqWuBNPydyU3tmoCkD
0qx2BtKpUGs2WwQ1ntbdPi3l7GCfNJam0QkCddZwII5ee9Rf07Thsks/MAjkfP8m1ZBtkNfh1gGb
4Xo5l9OPfP8n5K6AOKNgmvw/P6tByHKvKoOslq2MQZwlW1ig86+fSh0SQfmOdBB4fYhViCWxsh9P
+ZZHQMu1brBSHb2HCIXCMhCeBaegCu0j2Dh5RhFiHLdHUZ8FXRXbNUP4uCfdfcHprA5o6mcgO6eQ
oAcOBSYxoz7QbG3bHXHv6j8z8Khs68U9iPGgy3Bojn/AtgC6VmADXOPPzz0JaOjLUmAjWsU7fK4P
QaxFNsB2/ZvtxbQrqCuFg7eW+OwZq2tneRD7aJNiC/mlBlLzcdDUMpxv7UO3mZiLw9JOMwl+yD3+
a08/aAqcMMgL7X8YBmGQKUICLYxH4dORo/VFIGt4q0A7Pc+SRd8HGYvYEP7AbLk/DgyQhrwBzXsI
LtcH5YsZGykwDG8ie3oI4SBR5xo6Zj6YmxXHj4EuMEwfosW6fA50Pjn47y8a6eYnYgGN2/fiLstF
luY4Y4U44IDSrf32SG6JSqEa6yvIgYAKsdNcmLk1LlL0bOFxL58pThcz2fmJuCeRG7PEE3kjJkb8
eAUnCFWvz61LZ1tChIvlaM9B1himMaVliv5AhwG1tSvpfe+UyWaUor4Q8N+7N4mQ/XZ6Uf2rBZsV
4StFM0FXJTvcp6Nzp8IDCX95BTIM3ZsTd40haXrXGhs6UXCjcs2kuPT+Uq4ueEeC6rG2XGjutsXC
jK12blJX1yB9GGVCeDEveRaMcw1RDqI+jCblCk+oRn1KEELYDcNcLCXjle7kJ8uiRAiU1nLRp4w2
xK11a17TrWV56D6ML20tgJio0ALMG5msKBsXL18pfV2+1b0fK86YNC4aZOOJH2fS/o1t/qVJACSF
RlBK0woEzDEy0db9cy2vYcBlIrGh4Brh1cJdKC/yMduf3gq9xX2Cd+UGtjeESHG/w1Jch7mc4JoU
DUEfH6+mFn9Xa7xL81ET5IYAT5zyYpTOpMw4kytc0kjp8ujvX/3Kk6QJ/qIjNPnrvWz1eJ+0mY8R
HjgJegVFhADlYLgTe2kJMTC3rLq+VqOibMWXo7jx4sIGGyVjp7Mh0U07WVJb1AHLYpzNMVorhxtf
i3MNevWfSa+BS3Cvy30BJdI/OkhlUJdubuq+D55dn3l40ywhxcj5bNbh0plpOrXCuLFw4RQxS0PK
r5zFfQ4U5zB9GcYf4LcJKkMeegKwPzjjLRtI0eRMeJHp+GNrRtwfn7NlrJBQ/0NLipG2rPFg9/3n
7WKsS+LnFUvAoXmGNTQ0e1cMduMAIcPXC5oAm1CEiNTqM8MRxYjfSV1NU4FCpsCIqQhAiYYLSwfQ
ZZdSwn0YAWbYXcY31+itDI8e5euwt513z468xMCZO1aE0k2LMGjh0mGhfqMv7Z3Ysx/SOyGNIiNb
IMyOCAKHRHLpxuLHehyNk7mTbAil0Yf1gCINvKHDqJAyFqVJi4apBKWXwHmxuxM+mXl3fVr+rz+K
y3k6p/swk/iK+9fpb3wpTr9xdBg32eJxtfeJedl6fgiIrHtRNrnaxLLW3wfz7bFtvadS7RJ8gR5j
XCwXwerTDf4kMmtjXvquY1ztDqZGTJ/LD1gnkSyLf5iu5iJXdak4iEyeWmuoxWIY0Q8MoyUIdfUm
0F1uVWV3fxTQW2uN6ei6glf4khw0jq9kfzBslRlaRjaYkdd4b9/pCsCvLHdszRhqtVW2b4OSVWft
VSLUPGGwoobQEkwgsYvk7J/4FAPaJeSh2Xrw5iENpL8bRpoUTl+AtI+XNSMg6zsNWwZIrjQSIFWL
A21g0MOFb78C4joeFF1UL55s56uzEddvwnct6ds5LDyQYvwmVgQz3RG40VVuI9zPxu6f91ONwOJ3
YxUCD7KCFGxY1CL8yNW8a4hb6/rJ72cj5257lrHUaIT0JyRfGF9tW+rtnggNWNffKe9l4LRju5RT
Gf9gnwwOQ44mQRUBDcBYMH8DjtJ3oz93zNP3exLHvI1yEXE7iRObbqWJHP4Qjiv5LRg/lMqKv7J/
/cr3sqQjBCT2t6qq+fmQHJgqaXcZDQ1xyEYahmNBlv4l9n3oxV5HBzM/uZID94Pq0ze4XP5Yb/Lp
5GF78Qit+omGBFxs/hVeYPDhqmr0YzQtkh8/vcaE6CtcZuIoW5LfGQrvwuQDjHzt8WwsnuIAVfJ3
Xj3NlA1YTflyn6YjlJ6bfXEoZ7iRtrbiLvyKsl3kC2Tx++7ZVuFhF086CwuZfhjDpVU3VRh87ZBB
2JTlrCsRX2TvDyyTDIWJrPVMH+QctLTv4Nj7yj/GlaUxtFUERfpWfBH01PoyRvP9oKeBGx3pVL92
1qWrIuZpdC8knjzIuaIn0RBoTqLwG7gTX9skhhkm/7QE+rqdL8APKlJIW6DcEoL4WPCDzldocOCB
V9P1bnO/NwFK4AZh4hoha1oty3t4SlS2RxQthB7P7G0aYJ5RmJl4HBWmFJ5JwkR+K2ayu0BdmY9C
GTPaUzIXbIkehGAOj2s05u6IzbitXbmBnBDeMtRDNvg/eEzyTeXHdEguERs1kjFOUoEXYu3MWt+2
zEqgz1SJ2NIvEXz2pyVuvW157OhQQPSjb/Tw1ryl2JAL1pzO8kkDWBMiB12TX74DhmfAFtpewTVj
6ajR+KctV3/MFcqDaJ/Ld6j6Cvn3pptdkuazzE5M6FwHHVoWlc94L64/90xpGUMk3JttlvD/AIPS
HSmB8kufd5wQ6xrzJehsDZOngo1Cqqc5WLLgKZ6SRh4qtOpfgr5ZAHQ6idia4OzNEitVPL+2j7Wr
O+W8Jc5qO/EIidf3XLjiEXpjifvgMYsSsVyPjIZzL/AE9BCJ7+sn+xEtP5l+VTxx2NMPw4e1B0K3
0RQ/XS5vzDakEJXDmInwpIo6CWiB8fi9lhOWeTpTimvY5KWofs3du6DSKo5XLo8gIBxYnxgDh5OA
caWM0r2go4EllreRctn0J7Ys3jBCcs4Gt3mctU2lDE+7QGknklLBR+WS7idyiobvZCaaoZ3yNB2L
wxXn/Yb7ayo3lqkk5+PEBEexIX6xvzLLZGi3iDCgLVU9V0LS2ZzG74ssFOlLpy2f4AfAH328e0uB
qXD8DZfTFifLu1JWNR42wX+Mx81/OG98Wm1qkWI7VawtTxocbZJn+CIEUBOO1tnb0aF4qs63umlT
LOA/yy4tsZQmOYJqbuD96Ns2L4UitFEdkeGumJuAtU3Ba/kXQgh4jJFIiPibPjq0+e+7RGsl6lJ4
Kc5VrvOs14wDfZdFbOh4EmajD8SfP54iAeZ1PrOyX8WWzrsPxRzZwIJmqsC4zDT6HQO4tuVYXUNI
RjW/2ddKq4u7joVsUYV4AxV/U6LqQZjUbCSpi4FdBm8eJXU9KojJIENVRdhVlPy42Y1xCSSueQDk
7+1Tgx06Gt7aIGJMpaXQQjkTI8U7i4u+GDvYK3zbB9laSt88B9SvvlxZWmfbsS78ngyYaiilGsp0
gdqa13cP5KHtcn7a0FrtT2GBE+VkU7CA3Kv0mavSGumLas3yQ8/RKBhz9fKVOqNrEMpeX7v/3poh
bu0o3Kioey36K6Ol53+89+cEKFMyW52gYqDirVAn1/FXZUpe+gm3auWwxC98F7gTz6kNK2DsSLvS
IF8rfEHzCb3WqvNwXMkspbrfzYLOdICeZ2x0HxOYwMIDq4XpFZ5if+KsA4AZpCYzNjsJ9uEk3g1U
ivt1ajyx+5mN/YzcO8xyEIXl2nEFM9rF/z+3CSSpj/FsArXRVp4jsKL3oG2/mjdRuW2K8ulcLOPk
IeSvJWefPmvNbih59jQ0YYlX8rmULfAfoqgjWQh/CQ+2QXelMeYliavtTgT6vQeFNmCslRoyvNqD
2d3XsqqyzvJOGzym7H04aticGFpXmEFISt+BkYlzPd3+FjIxo1y4orZJe6VInYJq4MuFn2EuOj7W
IB1YPbVgXmFjaWliNXky5bGHGUyw/sX3ECBcYYeCCLMP/cCiBtaJk9RvnYG83beUcnM0zoMGHbo9
sDRCUFwvgVGu9jMdl1Cgvq8PFEJ41IMp8XVyelUeeApx6Jqcs/6fw/N5pDRutMqSV0L/mGRItcMu
I5GSnynZVhvTLM8+T7c0C9/g7uoHoys/THk6yerxTkTW7xTUCPvokHmD+Jhmv/y2zy6bguNPPf1K
i8QuBOcdgKQhVXVXAqqo2bDDdrOw/zBPugFLtLh2OuUYyF9aMQu1Ymzni0qOu3nf34od2dHMAEwk
3aytpeguIBHEdQ/6UWsLKz/eXTVVlFW16oNUSgYp3CPRmSbf3a4vs2tsEiFGxGpT9B+9rnRd/ltn
/kQ8GSkNVFqxHlMOaxqKjc0yChu/H9AQOpPa1fPt7Nx5B/zRoKBAganVZCijQRxXSRWb+YUoV0/m
WyZbL8n2/aSxbg6ZruMhgrXQojimol1pileqpWMDOHqJeA9bQ7KYSd/3S8KNkISuI+f3ni5ic+oa
HIPsIvfVGkBPHejY7ymNuHziDfCI1SDC11gM99Bd+J/Fsnv6gbfQrGgZM2oaVn/kG3nCw35kUmPy
PaJjwuTNPwyIMnklISCPiLKpC474L1gL5oeYSU4ArWxpAJ6eW1WSWe58Zkx4bUJPUKxe4jTwxj2j
E/1qTZFXnt/IJRto/wiLKqYmfkphUw/fMpxYE1ddDY2dNeJHYboP6GErBdf6Y+xDSILV2XDyNDrj
c9Ju7qpSlCYg1hZYiMzBmurJ7mqekUxvTBfhI/tfRnteaBLqSE7jKmIxTQoeWmtYQiE+pj3sfV1Q
6IUqulD+0yrOH1+59b+PFJ8npAgwHqh9/yCKLJE0jtpu0Pj0WtvXKNsG73ICOqNu/uXnglivoXr5
Iw4I3Mjn56ecikj5j0OyFw7wY8B9jcJgE6B7XRTBtBGj3sKjurxFPIjcraChrjCXtv1jwOoskYqh
ny9HgK1pAwHthsq9xW6mE7KlMZFjW+gpV9l0ejP3e4YbEUZ1Bh2wA15q5wc4xoLUOf0xaMxd2pni
6EKd8RW7s3fP70ga9m2InqAMCvnclXZUkY+OoLXuo0MQGPMGt+6i1isHkf48cOCOWpBuw4fIOT6p
VWd4BhK62yuKmjX0AWfCaYhC5c27Pbn3gOu2hODMYL4Lsuxk917zUJ9pFmb0XPVjFY/Rwva717cV
LF9rNXtkMZy0ni7bsbHhZgCJHoS1EJKhZztpBh7Ml5Bq7TGRHQDd3GEWbfOem2FDneUuUU3a9xNq
sXmVwk/3uDBqf3k/pkL9uEPjaG7atrFacKZmlnmTuUm7w1hDaF72yS5Bl2J8G08FXZo9vj+z8H2l
n78tZHFaE6N3kH4T8ksMg8qVoV3UiVaY7NtVBo46B0gZRPYBbCRWFRdhoufb1hEhUmzwE3F8OvLo
q99lEx4cxFq3ZZzYM5k6XO0c2My8AATQLYz0qCyL2GpHmdjPpLXIbngBqHMzy/hfHMdYa2a++R8V
hYjonFOrgw1dpy1CWhU2vH1l+xwhZncXACNR4NS7Zuat2gOv3+jQzeB+75hmwMZopbCfQVwK8Xdp
k4Chi/zZc0efi4KKVL2iC6+wrMT03XBIpK9+2HOOzlqbSDWOvi1anVJuagyOXsy44d0kiyCnmxXw
pdhwlJg3fL6VjKvJCpDqSL0pbj356eErsXdn8SL2Jwjctk8FgxuI0JkuBWDS88GDnus+xzBEKgCW
v3fVjzMQluFNyjObmECEDpRyiHgolLLy3X9dR0JXmv9WmyCgBSscXeNaWBjWKQn1jnzvOJ8PTfO4
jaSLWMKlhl351o2JZXhTAdylr8Hr/Nbnxnqnhs4NLOLmZzQBzcu/xSX/IBLLhu1u8gewABkQpDgQ
wtuqHS1SPqZpRqv7TeqmM8FcSvI3A38Sm3cxTO/F5qxR6xcfgs3BWptDrPr9EllOVMEaVKt6qMlk
tlhbsv6uqTXwEehUEs5Pk3Wc5unkhekHkQIQYG8fiEsjfsJGm+rsyxVx+v1BqZWU1gHREiXqB+Kk
eG1yx8dwjKg0WXi/RLxB5GcQCLYzgIuP7FZHQyFmv+UenlEWRWGxZQw75RTv30f/I3phIQsh2QVB
o/nrO86tl2A0Gqkpmux6KQp6hNwlb0lMT2ZnKS/GZ8wLAKMtc9NET0BOi9uThWwMEVHBg1j/3r1S
0nyUYb6m9r2TBtCFOD6Gz6bmT6LDXkmLZQTeT8y8AeT+pkz3GfyMqyF6i3dS3P4RW0nC18IXUokN
UUC+V0NWpvQWVXxDByepYRBdDtNWAf6NfuX3VDpYUWlLjO5W1Fgd2Ip+NIhA/oh+w4rxmy9kOn+S
P9WsiN4iIpu0CoQOh/emLUkJfwAnYZnlQf63eCtzhs/hbgT5vy5bDEVGEpgTpsoBC8yeu0nc2NTT
QZq2uInGAqzh0UozQrVsFFk+W2/pNl3dTkrtWeqT1pbIrRv1ijeNwKyJoGWD9wHAvuvVEllZKvr4
odmI2Z2k2InaVE3Vg9WogEmTistrmtKaSL1NP4qHuh+rdW5LFtQv8WcWS3uJN1dfHDEiG0k4utQh
z7Y4Dqred4kZ8pZngR8kvmBcqTFTydFp1Vqsvq9E2mWnPGuFRu13QY7ClCNdsXgsDJs17AjE4906
0MulYk5X2uSEEkDUqPMVMPSezU/TxOgURV99Ek1Inw3OLnfm+LLyXZmPGaw5ZTyBdoO+fYZzcTOF
beLZ32oRAz8S7fiv5Z06DOVrb5jBF8Wf4lcAfmAmAFNuflMB4GxnmVBWLMKTBYxsykUbwx8wL8sf
/ZrBolRsgvTOjibqj4HAnIdZh5+8jzBMeFCWZst3tdKrrpYW/jEWDaUrQ7WiXmstitDyB6e5qA2+
sZPneX/ywPQXFEx+HCWA9Uu0H2yieKQBnN3vlpAtY3ekhae/9Qi4MA1pvybxHIvbmQFhfGsOTURB
28VgPFdMgJL1+pKZlIM6qROkEl9ZKhVu9+UJkIJwVIW+rcLTwwKA12AnBhsrsdsXskWduvj2xRb6
k2hEGucTOvGcueYp/gld0u0BEm9f/9mQ/5yNMCI3h598T82wD3YUkXFHIGy66damsPUhOLaIyrqy
ZZBy0fEyPP2yiopNHVs/hZl4u3CWGbsJ4K8Shg+K239IQLLdGS6XyGhkieweSehEkZ9kvPKDpEWy
deuYulVZ7yO2oq6+GxgBPk79uq9NuFMerUc94sMzJv3WZhugmfG+UuEGOBxtpQwUUcZN39QJdx5j
VIPfY33SA4kq8XOIrWXHKJ9rsWuGwzfyPHD8MlnPezNzdp1zVzh60iPacDXwsYk4sAs/RsyG48xR
qewVRjTuovEPstQKLrT+2gS7XCjB0UeO+yzbgpLvibE901e2IwmBKNTDwlsej30nsvXQAw2IC2mu
BLoZhQXFBhzmeEHCjmRf9tuHT1ZyCKHB8g9tLJyZxUUF2yWl1QsN8VHPDP9E9Oc+Wb0bHDrc+/2j
LvAkZkn7bwLFTnwfr4O9X83pfR2ePK68nCkHtRDrRvKDUvvzwjJ28CyQILsfknt++IkSUBnNBwki
T0jY0VqyxSezmDJueSuN4+th6+kXERFneYYfJ9QDLVGxGF9HuPxwj+YAz9tM375OeiRpssAXqROK
trsTHfq5025S9pBkfv9qcwq5HY9gWdKfzH5jVJ1LsiQUpe5gQCuS3KClNyWVjfQZJhwL2DG2lnjp
/apWpm/z13Lxj2IaggaqIBP3pNWrhvcn5PJKc/xzhi5J707yZIeKW5VHUEyjMvwvrInHx21lRfwQ
rnbE/2SzGET/uU2uhQhI6dXKIZartt+8S/IBOjhG/p9yE+Ksv5oVGHPAGbV1zx6o39z+U7c2zbri
oyzSjjFNxDwUxaRrvnXaUQ/jp5BhjmsDTm3/bDXkzMfs+tegja5Ab6l1W+ateQjDRMzh6vq0u2ij
AxxEshlCh870ewXwOFUp+bKm444iYDr09WKcyhpSQnd/xok24e26t12BE28mBNMU+LMrUJFmP+0S
AFLnl/uGNt7KyZfX0+B3Ir2TQ0EJ5v0SHW1O60mClkxEBitc08rBM/N+GufUNCAoNEPfDv7BtXGS
lDmh7FL5spCprMGSgWG5TeX1WSmEvBw9uoS4COZj1sUuLnlWEwX7vKdlgNuBofSVzSDNxjZtoK0c
D0rkXI/Lk/Ly6LytfiD80Xt/RDscH8C5idHvvWDX3juL5grRocNvCWBUyNvwv1StPQ9Oz8LzgTnu
EtCMLDrF7+nhuD75vzKaRrLcuQgmBxPxa+wQ+EZoBoXDzompT5eVczgFerY7vtZVlBxdTWKhCJac
XXZb3eFyR19YLb8TsJnQya3c8cBHkP6JExov2CGrlrHv3O/hLikO8zg9zTu05JJFg1/PkQ6BpfvF
EkRQfDGO2o/A1R5QiWnrxxtnny1ENMJ/G39HArUaQMlf9TY4DJ+qxqg5JSzm38VCvXo40ORJyiie
u3JPnIYgz5T3GZ6YktUGqeJUqPqM49accAUfG0sQAkiyTgd5eWgcivegcZH6yoSK0xodB1s9hf0g
q8tjyMnMAPis95IbSPI56eoYcJyf/oXX2BXVUdmo9ECc5aMjKHUnPLselCZUO3yO2YoJf4LkCuJL
16vhsW9oxBfw7QOVE+gyfDXlSdp8ffap4PO899kElLeSlAdlVko9uuQc4LXBBqdXcXpM9eLPUYVl
+vMIwHtTI9MG1QP+SUtiO6+DJJQJLquMCmniBYVmeOc/ipfhmqfBPm2KhOpfAjOqLAhXcmP5BjDB
cZtF02hg4q8m9ZThmYxJHVC3XJ0XMk+2hUY+45EyScEtOHI8pni0I4gLa10tT84jdUhsFjNZAgSk
1Alcpgl471dsMq5uKWyXAovK7IjeL+VqMjOcTFFDymlUhF9pLsYApPRUicTX+Gn+jWOPmzAn48Pw
FozkPQKZMZsxhRMPJsrqenNysE8HY2Y/R7MUUgbs4O1kuq/d6qO+nes4kc6qkLjfCnQbz4xE1w0T
+4coNS3JateUYSE5X1I5sO7eNH1J5mALxjj0VPnPicQcgM8cUW9s0ql1NayuxnDxgPAZXL6bW9SE
JrquBRZmNVCZduIZkJXmPtMQX2eqnVCRf/DakNGqiQr3oOn3onfyYp4J1QM6dI4k7dH2Flk3eZtd
cyDoWrWHxrnYN/CECjIjXxgkYVe6Tq+2Euk4dMbeOR9JCNA9h6s0AS5Zlz/19ju6AhMyiUIzU+BK
Sa0pK11+pJ1FLErzQvE+YXqpxEqC/6rgzMt8CvyuPxSBnM3Hs449AbbPBdZ7iFb3GV9PZk+zTwEz
OL1GUDOC0JH1iZHWEJZQ9lNbXngz766paDkhVn8tKwXG165ccHN6oZ88IjBgotfjSoO0feMB5kTL
X2wfHsVJNyPxxKXCWoJYXNnaM4RpUgfhy/eahcrml1ApFkfzT7Xql68SN0neSkptTFkhBS2OXO3e
leoZcsKn7vgoFcaPvvD3gKxspHzq5Ey0d83vOR59wrvPn547/V+waxJ/NagRmdunNbL+ik8lwrCA
YdAd6uGQ3bq1f6rFcpaAgH+wll698Lo7Lcm2Qutla4emRa6dCO62erGeYp/iAsb4pSW2r2FusL3o
vcaRmKJQ/9d3RLS/89B4bFA0jcrS6LgrehKecHHwteZvOkIhMFmNy22OG66lN+8BdWNUWXgPXcgS
RzWe40huEjPkoG7XnPKr4OTz26fBktvs+jhL5VhNNmYtXd8AmTFjjLH6Kum0kA6VnJIP7Au3jMLO
ncNa9H2WJr7kvqtpcCxESbDAym1xXpvc+ppZpXkYq+Kqvj6gnPGHYxYod6bRPaUqK1qSs6TRFGL/
QmGfYVSiuqZEVBorGjitROb1SY2Mt6iaLfhLicmjcAG5jrNBuKFTm54Um+8LdNI825sS2A8ch/td
6VbRLpFnuDXOUIM7F5XHWr0/OxLUNWvBxeAdG9f+iZZZaUn5Ul6J1AWt7icwtCv5x4TRNAALcQ7D
J7lHuUF/HxJPb4gNolwzW6KGffu8MyV87ByMis/2HxxrVslL7rUo/jD0eq6xkXaisiUBZdjDPnvR
L1+Loc7fkBlZpeQmGSUGI/PGSTVvYBDiqwCTuinmjTjbhmR7AnribA/lBKlfwciMMyjjjUuY0JCJ
p5tgQMXYq7OsMH4C4rJS2MkFH4pejPUi1SJh8ldLi08dJn21kkRNHvQgeLcEM8gASxHKuAzwyfZ0
M9Q2kkYJvC+v/11tvJtV1JtC4ayuCzXDx2WGl2AMWEoDIEIwD9nq1qGpel8x6RDI/LkkrgTq6Ur6
sfQabbLZwi2WK9bEI7P1WfB6TvhwCMJH8FHPqjasGzidQTu1emrHV9TAzi7V0xeEi+d1sB8VlBrR
wQEWUG2CWRTF0JAH5OWwxOkjXRMMC2vQRDBA/Qqd3nByysQn6HKCyx15RATQN0Ymq00n71Vz7p9o
FteXD1/Ikn5W6rJyL2nNMjuWjGougKhZn+xs9j6SjqK/fMMQC1K8IJHvCYkR67W6u5Pk/QqfgwJ6
p4XNibSqyX/MknIYP71n7WICt5jyoqHb1VJxEitxYnAgSgcAuaK+46bL44OsdQrHyus9/Qxy/u5s
btcGGN5WjCff9zGHQ84Zi+2fSmZTB3UPSh+uw06mfi6mk3FtO1+vhOLdfnPRObDcDawu0aza74me
G4RnR+GUYMOE8vRgGCiDJeNMVRnC5xAJHI0q9TscbaIC5RM19smDRsup5dCv/CVxdp8wP7cBf3cl
SrCuPJ/WNUafDOiWWAycieVWcS16IUL36Qa/xQYmsYxeWZm0cs6NfGaIQq1qXFkB6MALoeB7ySFJ
nRzbP4jNO7bOuAoIhaHwz9gCcubLqua37Bk2l+ebNi/jiH6dCwD3+9DQvGHzvdvEUBrDoC+zzX9y
a1ba4Sv2TaGADkV4cwmu4xqSYsPJPayGNYk48dcoxHDlUO/+58hL7NqUMTe95IphqV2WXnWbA0Ik
sWxsCe5I03OtVUsPfJZjnTYgefe7YfgepxvFZ5fa2vQ9DEq2ZGnczkeLsKLOnIxMEswWn/NksGy+
5dJ5W8ABx2h2+aT9dyiuZWPjTtyNjHlqN4gEa3OA4zO2OgMZ9DQUNrW3uKfES7VAdSB6Iprr0tQe
ii+SR/ZzcqBsOtWybC0d8WrsQgCyNQS6RpbgSzT/oaHzuTCIl0i1mrHm2BvZ6m5/ymRM8J7IUN0v
iIB8Jnw4yGdOOgPyrDVvUpX3BQYAx1HW/JoUIBNHnQXegXDzPZc8AAnIRdiya8mU+b8vnf1I1+et
NrM+XPf7bMOH+0MBv3MMebyc1auTkAtybDfWmdD+aWkas9DrLUxoD3dHgZat9ue0SStRiTRCTg4L
Vw1NB7gX86RapjDlQZZEkFOjYcToNmqrDjD4sAapKrZ0IOiJ2IFfTKxNNkEftos16kxEBkXalwk7
3yZ2l+rl5g61ulwvbiEKs97eVpbF0BUaoYN5ZJ7dNV+k0lm/aARgFnl1xmKX4jEwKLzJq5z4Fmz2
7w6Cy5PR3/OFLtURBvZ32Sl90f3LzcMFkuhjjNp0G7hDCe2RutD19B2EbV5JiZUraKZcZAXZOfhU
rN/Vny8KmPgPGxuPV2jr3l6Mm1qZmwGw16wK3tKPFu7vPWWR3Dfhg8NQnis5pvLRNASQG4OaWtnp
QvtGDBVRiRCLkQ+W04AAVqINt4Syaxv5dLfJSdNrGxU5POBjUK9dBGtxxsj6meNL3TNLc1u/PHWC
UmY8REfL6AN0ruFG/ZG32BtCh9v1kc8kxel+5iT/0to4AqSByp1AC+cjCUauF99ixXHKYCGwa2Ou
WqyCweMQVg+F3RvoCbL6NXzuHvZ9IE/1UG7Sf31+qGos/CsEcJh/3ArKG2XLzoyOQtNU2e3/Qgh4
V/3SU/ZwarpyXZ9kLfWzpwhy+wRgQ5jBFd3+Qgjur8IAOIn0mYFh+WEN62AaUswto/szwEvlRcMH
7gTfaQAKqPkWhK2Wra81VcdZrIeXU31s83WFbw3SG+ZCkhuyWiuw2d+CGf33+C9hT6bzkODQojXK
qYFJf5nmfGuIYxaqJAqkqnjLTupx19TYunfDqspWywjuCJE8zWQzxekzWwzM6PiTDn80BhA56/IH
ufjerBGmB6qEy9TG2joo0QqqGTcVdJ0UJBWVeaLR5M9Egtkt5bJ9PYZzCf47Fqzx8fdi7dOOfd53
i9J88s2WkdsVFxBF7/QCodW1XJUVgZ0I3DYQxHVKoTCBlx8d/I/RSm5zlr/DS2qLBsgiM84GWOJf
bLoUyQkMXp6D7gv3WQqxVTAgpymdCFX0M661zM0xffUldC9AI0CMY7w6Nq6HCNq7HY31eJ2gM7g8
cCpe1BN3k4Ehr2FwlzrSPK2jD8ibC1BSLpgWMYw3Quw9PYXEO4zwUpM0L45SHoh0Uj8J5sCdjqJB
3F7UOif6RQyxOF8ERCoebdlfB70cAaaQpnIJ61CY8fkMGPMfDz+aRC/Fg2WeV1MhA7mh8n0zqAmP
V1PoEL0Hfb9+OAxO03AhuwB5pvewWC1dk0d0UBWbFGFElwPUeDSlr2XLqrjcXZ2QYZB6yDMJ1pSg
iAAwQrFfSNBLbaC9oLgHoUsnuh+0AeWWwmkXaR5LWpzvC2S4SjZBC889QTyX4W4lHFJFevU6iGiY
EmFzb6CIGIfInPflfEHb14rQdmaFsKtAbknZYvLOVydUmio8k/RRNlnvix4oC1zpx+OAKlmosblD
CaydBoUauodkvQhSXccC6Tx3WL+z0U2o4iKTiHjEjkhCkYHDmH+e04oajUGRyL9ihoq658FQIlQo
xrjfCYlBoklnyiFL85RoHHjfjEvDeyoGIxBHW7dJPOiyQ1n9sf82YWgVHP7pgSorZO9BL5rwlltN
0aOovkv39rHtmQ9AVKLhTdxUxxGAKPeglPpWDMPh0K1AAHGwAjL4HBr3cH3brvbe97Sx6S/qwsqV
g/8Q470hAJHb1Z9O/2bwYHiV+LH+evpVnWD7uWQj6zj0PMepLJgUb1++bbDFmSXMT+Xpm5RFXbz4
GYYRbl0QqgYG7PRCVv9gJHhCSmFpmv/WH58Aijh7k7QfIpGAmv4SwcRaDEw+HM4gedT913yZzUi+
7GE5xg3tEl6fVCvpjfoYF9gkozKtub0YM75FwCiX8i5OYvptcwMN3U31+zMKCUow1mLv1nejvsZY
E5r/LOLwhr1MBvHGu+Gbl2SERzQNRMTXdeIxUeU1QZYMpwS+zLobIs+45dJSUpnnlwYNvabG6+OQ
IhqlaY8ab32/VLdQ/0qtIC4Cn+zZIQHrDYyXddhokK0Cci9N/JmiEHShKMv0joCz0bd7vVTLUT/0
JSyekAt2IKSGdcG05EWOXLJeMvVu6WOfd1w3vTBw35VBU4ETEE55tCSK+1QPpeEvWUDXvKoVLIdO
2i/wgsp2F1Bx6Gbw9RR6iUbwNDp4bh4pWDU6sF2ahWZuBOpXXyV6D0o4k+J09zRHu9XREvd/P6fQ
SkIHBALwKzrdeqWRuU6KsfI3Et7DpCgcnOw2/NkMqn5qSW6une/2KbUf/omxJG9yR76CAkmQleLi
cQ6P6VhaX+sNB2ulP62FQ7MfWGv2vM4EdPouNZ7VnVtgGqLbwpXYoPgzyZ9LB1ix2WMv2mhDz5Ib
/cjwt13ay0XVn70RKxhXFCvGx+K7j52YISDokWEwwt0AYg4a40lqusxV7a0N+FdRosNYYbUasVgT
G1nBJSP2PGEo0B61lTz6sYuU6sg/PEM50mcOYDLqy53C49SbE64UuzbsiSYqoz6bkPnLuuUShtZR
6faKFzNsdu0U5pj3T0gNtA7LyEz3fOiaAm0H/DkIj9GAY0jRPvIdNzgFMRAsQV6pndl30ChAgD98
V/URjEVUyXHuKm8kOX/9PTq/dSETwPgNIaq/7Lk4yqxICovzEXtzUYaoqmLjPmcd7EGHGMbsgXjM
Vx//tHAU2BmHZumqktguqXRhsZ5t5tiL5NbOAAD6FeAEq8WASgwkDkF/tfRn+1/3gPv0KQHDYGOb
wjw7c4AOJkUiAHxd62x1eJ/LnYT/S1f7xPZfjfP4+w6147fZZlIOzIxTdKHv/9DUIkYnoTtjCSHU
8kIHjHS5RoZqE5RN27zfRcK8G3XpO4IuJoLCAXWneSIeW5RW6ddq6oXNefzw3gc1FKh3ODlXRpk2
roRnHiMo39WEa6CeqQPUyuKmbBbC73Z9vZVruMyPczMdlBRr9scvWNFPf1SDmYPio3tMv/MHqxCa
ththsnEkIE7U0tszk3nO/jfQz907RPAln13xX9fLU4U9q8UuxR0Zra3JQrZdOMXgqqdtRs++wryP
Cy2dVc4ap4t5pYaT2yrT+C0afl32pOtUUO8Yya9wgTNGH3HmhRSRZ4sbRVAzztq0sTJ/mJhDC9RA
Geg/lnk6kM4OekiajMsyNbAgIOAnDvVNQGasluxsBTTuaS6HtFRY1U5b1P/IlZfH0luq4bDl6ZdR
j2XcWlcw22O1rLA9cXJQd2AOkuidLMiNuK7IJiq+I+2h/G/UWh3vWMS7Zf5eRu8qnQpMiz43DHC1
g+q3oKFTuVkKJR67eYyfwHukgg8dLDDZgAlJCLfBdRFr8tK7Afq4xQUQLa5XHsMOQ2puMAumlpkm
jMrfjLnvqmMwyJa43QvLFJyC2bXPnFbx9sIf+3mffFi9hWgWlF/MIwF5/+odrYKr02zONP8tD+K6
9EQKagrekn5wgxWN77LcXwdt9e1+vqd4EtoPhVfuRN8zVSDieoQroK+b7yvcx+XX23irXbBcCwKi
opes+DvpFCdTR8di/Vps6GwmLZ9DObEdRSykWyx0PUPBIxOTXwgoQsAQuvHACXvsdP/JBjvvWkln
MSpyS3vxtE9iPthfTexz/FAwgUDjQSNonteFg+vyoDSDZtRXDglo7AZQ/U+if+Cgnqk7uthIqsNW
bywcBC2x+rBbmyawv/T43t8WrYx+5qf0OjrZf/aB973lQCxP8Lq3bjeVIwdSjbR96o9tM8Bwsw6E
415tCitMvyjy6oFMMtmCFGvs9+VDZi1nI0tXLE+oU0MFnFzqibXeoj6kSUolXRrA6cEGRXgaX2uL
KEEtt5IFgbh7h6YVqcvXOBgGdtGqYrWKowlbLZaiuFPJs+pntkDPFpLXWucBlUwxryaxILmxN1xv
SmYCTsU/6cjCwZ5fCSq2xv5dTxLlhx4DuF338+mgBVI2NEmO8nKxTux29jgolwI1sqApvX0/y7AV
N9JdNuZcP6Vq0P7bs7fvYc0uaYhzuW7uxrPy0cAE/KjYWy3YotN6aLG4koAXeLVMyHRTp2W7pTxp
lYW4BQSWX1ro6Gj8qZIAvn5LY0PEEHgDbNyCesFBUeJeI8LByG235IKbQmmLyMsX8yaiaYLMj++5
Shgi2BiuksAkt5z4+N90qfP8RdGhh46fSF+oyo4LcK9AejUatHPr5iDYAym6BTKWms81uVfr7nfz
yhU5FvZiQckPQLKSApGmaWj+gPRqz1c9En3UahwsLVXjJ7WpnFGY2C9QfQU/RjuBamM9LQGLeV3A
ytCbSpnS72MCdVQYaxOW2flwzqqa+S/kHzalb7TPWxNQCn8nEfuOD0VHYE+8I6ya0L+w9DH93k/q
ncHmg3OWDUUEFrUSLLBPQtcvc9YdpiacShdG+r94ZpvI5JjAM5ijvtpL+4j0beLl7kjRF+E0CUYz
Ud40WDYlfC6TYHWRDC4vrnekyLVuNv+sQaTHcbnUe0T+3tITgN//gRee7Byw4A+QFV58c3V0RLJZ
RPKJuzk0klWh7TPt7A5NH+DfuWp37u+ITJFCfMoiszg3WUTPzYCMoBr8sLtss82V3yDgCYa9lHRL
9IX9xSvqUo9XIbOVNiP+BhRRzdMFoe5+rsnOeIzs905fxqywfB8nmgf93kEOCjqzt7C/KSn+ghZE
tFOx60beGBt87dc5zlWinSILYigahy20jwORexvCBd2dJLrkj8otMX3M3fmwhxyj1DUQnhskvA7c
0SwUXNpdMity2OlhcMtmJyKxs0jb7aT0SFsi3npgYwEjb1e1I+8YB+JF07d4e59Xb66coVTEAfGf
Ai7ezd6doSFPWyPT39Y/gF5FP/WKz9z81WVHYYbWYD1p6nvL8I5YD/fMjRPRzyPX1vQRnMR/Vd5c
5sZvYEyvjRbgV7rbCTEZ//ZVIXRw2BtcegwNgIiOwVsycdMN/OaRE1c3NlC7+DZBmiVgZaiWbzK4
WFA72nIpioavLvealhWn4NRmeZ0uBl+sNzy8dJKLTU5EGzy+2M8/W1EV4ygTFob81ukieZrvsIbY
Q1JGNeY47S2pW3i8cyNtaioYfCDG47II2MZu5TQ5C6DNyzaOI7im1a1LjCBuhIYFn64Lm9/3RKd+
itW310y5vG3ixUgpds0w5qf6RwAxWJho0Ig3/vNWyYI6ppRXumY78D3lGxZQ9quvmH+sM7xZ+so1
B1geDnuilWm6t1WoEAgrEkbCRhPJLwVI2ARlcbTGNlAShHqMFNalbh3htaoUCz1dHRJnsqupy7oM
K6FfJEgSIm9WlC3q93T7Tpuvsje9+3X2dH5yRxutAxdmGtQ2uBQ2gPXnpv4Nx1mBwyVuVbAQtqUa
qIegHPHQU6H1Kb61yY+IknSfhUN5oS9ouD9qREyV6WuDDacwMaJQzn4qb+6aVILU9fRfP7ygP0n0
crS5FBAyI8V2dQp9Lf4pThz+kcM2CMCwjeRDa0jUd2KIUTup5yZyQLL95LvwR9mbU2vnJ50xGBHp
T2QqBzKKAf5isEhL0eZ9b8V5UvTyqEZ0+vGacs+XsYSO/ZccqKmvF+3vKqgnpTHA0LMxv7dXwLAK
12q/l9PIkKwkNLjUhWY5Of79HlD3osHh0iy5X+Mnvg4PmR9p/ghboDAdLV0ty5pOCAYgLsXv/v2W
KmXGndJ5c3YGedB3T/gk8pXxmVCLJRGspl4GkmUHS6yefpWiSX+5Hna0rAiFGWjJlmjPu+rtBgk1
UQM9wlMpRCNHD2NlX/Mav9qQwqZfl5wN9NGlu+IttAFTDc/zxKeLRaO/JRLbLkAb6mI4M7aOrNnA
7wTbWwjJJKOeEernnzrw1Dxobc7jwpjmuvT49o74hrTO4Y4W1rpOYGh3v0GosC5M9SU+23k69AiM
CCQYd8vX7JPGfgM2Fa/OAZ5sctgpVPoGlW/FD8P+t1pXQoIAquxV3HrncSlKfzhgflfmcajc6+0e
Wa+rkD65tbo8I88PERUtK3RKxIH0YdUCzc+ryIVXDA+sQ/0lc2j17x21fHK1otTT9Wq8EbtcYg8H
1ldO3nLXs54PRBx/H+IHUl2TcpVrG6Nyuzju3RKuprHIiiOYrWis9BDL/t6XmEqztcATf7dAtGS9
5iHLZvwKmUpqGTiS/VoqocAtmHF4lCs6h09i6v0xjiCzxBlvItXLdNXaTt4qmrvoAGglaV+KkKU5
xS+WRgpOHxdPtbEHUjkARsLiSTUA72c3kbJxI8uaf5g+Em2gQgFUgbtWCCmrAZoXjvhqiKCaBzkr
k0z/ApeYZVmeD2cN1D3Z+hTeOGBWJMz/Ifaeyi8oV6sp/2Grs3Da3PEjV5ujNTqU8cWz2xxMoeCi
Wj54WO91fV3W8bLv8/vEhnoZdOj1FzcFVP+507VQGMNjdr3W/ejUNS7KPBTNF0kyo6zspUXbzC2j
S1K+jNlHS3s4mD1obbRXs+3PTN5de4HsXqK8FVwAWVkj2HxTJLxAiKljAW05fSFP/jxvctghg0W/
S6IB2GMKMxAf+UhflAxSke/xXfetxNMjemI8vAwRAJFYdZQAKRiSGwuPgKTMpHMcci+ZLrmGajMn
yZweTSTVLv8Qswmanptwfm8hycoFN8jMUeI/0jhGZb4NDf8M7LkOg9H3tgBGyoLmqu2NRZTCKOJo
7ghqfUP8zmEs8URqUnNOO/KdzqocwLNMcQtus4CxL0Xt7M2PD0s7QCckS8yiNTxrjwlZLXkGKlu8
9TBGOqzDXBJ3v/lcGqel/Rm2BqjdIYNlL5yFyl7JXpcekIbdzMVwLZn330Y8g09/HLuez8qrsCgJ
vmubmW91152wq04iaUBXyBWy/fJcufRrnE2nVPr+E/9uaa5ootOJp8erKVKQb/clFRQuWRfZnxn8
bEFsG39Oq+tsjAci0HXeKydLXw30KXpZEK06wVq7NfrqPaARx4mLWRF+Q2Zfzk6ypHW+EOBvHf50
mbQDiCGrK297OGMAYAE9zWz5MDFvIp9p9fyEYrTYs1tIyYyCdAY5f6LH1KwqHE/iJkB4SpTUl1iW
Tra80nAxrLq/VY8aFHgJ/x667sgQCJpUPNv9+0NOuKvEd/gl++zjAeZgUVNlHDaiiQ/BAjKUjcnX
Y70/SEiKbQrMGgBrOlYW+hw1E5Ei23Lk+WW+A0KiJPEFtcQ2EC2TOMx3tdxoSPGOeg2OL0yI3XqJ
LKHr4vK6rUXnggYyODxs5sYPaY0DG6lTbumXzKzjEFZ/Oki/BOHDtRP4hM8DaIw9/yF5MjHadolG
QsvlpVWaXHWNDcamClTBbKMAiwaWVBs6rwHbdijMT3kaH/A0LSmkItyrEWTSYJEPWCtdqd9Rbbx5
jUfyAL9b8oncWFc9wtvg7N9U/Saa8VFzC99sK5mSyqsLoXcpnifaNiR27B3ZASVuxxPCeb9aWnBe
nFgQ36zNfCRBDeMSxNxn3kmmEZwTtSKvMWslbTTW4Lf1N2dg9NL+8jJy0WajZJqCGxaV8tC2OhP8
VOYfgxOf61IpJ3p14WoKc4MJnaaR/aVQaaXjXm2vR30Gt9ZHsoijA1ljjsUhfGM9Bn6Pc1j55/fk
y3Q+v1aWiaHUn2WNAPJOWZIr3GL0iteGjT9f6VDnOQRSXZbntxmVIxlJN6xR3PjSymwOWpQvz09R
WDJ6wsAlRUD3HpPTQyp4SECyCZ/oMgJhsdd6Lv2wVRLrZQpKAjCdOoLlMrFAc6ZqCPUyIlZuhD7D
HIu7MMDjoOBwX/YJa+naEKrQ+9OBcGwZSZ3XU7hHzZQyzltvHfuu656N3G7mhbPf9bb6OoCMJxnh
L6iZETNvTfQbmRmtQ3fv3O/az992a/YPImVeiwNCymRvaXlc8wIZH7idqwKpDIgvv7crdm1RbIQW
cwpuTtvl5E8b8CFFtTr/0kGKyaJ0rAtgj2oV57qyWZSnIfdsHb17cCG3pEoTp1FBAc4A6eu6NhMm
PQ3WVNyfq5nmfkGTO6hOHc3WT0PTO5evnoJxg0yosZDYpZ1NUNbIH9wIGsr91x5lKLYrJveXhNLO
ya1HQAT8oT5XT/ebT5I5tRY3duu2gY2W2R1a/kwNCcy6+PDlJBgJvna7BUJf2a0uvOuq8AnwI8sB
fpe4kVFArEwXaqOSVxscNc+96YxemahDcVZK3NlMBoymFlxWeo0H2Twl2DzYHkkM7L/G7SPJr8Cm
GCStAXj7/GQNRBCkctLja2yFXk7qZi/28+6VxIBTrxfHvKc3DaxTu7zNfww1kzJ+Z6WenEBf+46d
DMGKgfyq4bhCYnw/4X03t9nvR9wh8qw1jyce1Xhg+7xGlhiitAzyPcrsL1EqE5EYcRA7tF6JaJqd
5fbjtI5ClRVyBbBKAhy0dqO7/kt29Y3ypNqwaoVaQUKDsTlIbJwVtv+P3B5mFoLyCEnqA8UsmuoB
HwZJg9VZYarT49mpfkQw1VCF8RP9hpv4211v6DBaeU/cODjDZ9GVG0OZy7sfJ/HQ+/6/l48Faw5f
onrdWlFl05qHN0OokaODq0ZrZ96Dbp2xHCxmWFohEOQCWdcFrCdn91QB/lqO8ICLRDbG3S6VnvGX
hFjHKzat8M2u/Cv0gzBsxzlr2qc7mnHj5OuCa/hAIb035IxchxukmUKCj2xukSle/0WTgcXDDclJ
s5bW+PDAAPP6GxH5IIC0db+mfZmVYyz8c+fcyf9zX0NMHsZ1j73hcKGRI2lO6PBFnZxOFObU3WHm
1QSNh+dnasRu9OdA/9qy44+sgHHAxRBljr8Xmt23O7MCBBAEdNXNcvMDQ7eOZY4c63JC5SDyua2i
RzQ/zRwZT/rJvg42KiUQcQMQbz31Gl1sAD33y3RcDsKJS0WR8yZ8BNu2FIgMR5MJ1pzZ0RdTjwTI
hDJOKYkouFHvoqDVLuZVmvxVIkg3ih7a78PrNgsapEtwCF2kSWuaHZSJCHpc/AuT7jj5ZKIqrFDR
KJC1ikyM77U+pvpWqiQrRWV6Wx2FkL6jkkSixZ6chWfzI47nO+4c7yI1UGjMPy0QJjnM7AgwijLU
6+9cSoiPhvzcT8yMiNWGC01KdonTCsePUn8uwFwW6XO38V3+uYXR42q6youX3AvOYkY1Ay6dVXjW
rAqK8FKVm2zoZk5/I61Azg/QhuFAcpNd7n8720d+Sd8ua/JhEpbSZsAYn9ZPERt0jr03Ve4I7TU1
dE5rrLaTeNY9F/3tCrho3YTjQponl0GFX6fYnassEVjGaHb4HcNSddYfPhbswqPmD+OCvQf5D+af
4mgAgc6C0vRS5UcWIubpf9eLixt7mcBWbiNFBI7QmTG0UzEkvat+Lja8sIqotTQ7rwGl9HIgVw0M
gsxUyCdgST8q0wFiT4YSa3inhkxeEAhVh1rI/nw5PxtbgrO9xrpmGQegZ0PVlXgUaRf+8gJpjuqI
kVQ0tUc2UgPhXYfGmgOK7KldWI6GZPeZie5FNRuT6DuFWP8ioYvbQHionM1Qat83arLmH+zRE9yO
zlHl45k+teCMNqIxfQXgKiGWhhiUdeTEru67+GAShRFqBvb0x5s5aEJUHDNsdkXfj5LbH3xE8nH7
j8w/pwDrJ5+tU6soGtRvJcDuiYh7HdmO31izLJ35Ed2QFEZHae5ZF10GuILqBw+uj0UH4p55mlNk
y39Ray4ax50Cc+zQ71GNuKmYA1WdAhxFNOczeD/du+kTdaViXlikgJcVVUVK11hnh7XL+4y38TFK
fDIpNiyNaAcblXCa5zK8X1kWDGxOQcFNpBINzaat13kBciHCzU4McKwi/roRpIrAnIvW1sGLNdth
aPxm+UvzlKT4NYOX1afwTZTyc5ijs6bti0n0GFb0Mdos2N3YP6dwywmVbRsChGZQtTCzxMFI9JR+
35Y6v3TAG0aTqNZ2c97RQVIXsMvSKte/TZq9IwvRCyBQJ8Lo8QX8gkwcoj+AjOib+gIUdAU3fSDS
MAvHyFFxsi699x5Vlvr/nL3EEPLxBq2/YaQsxTbNsjcBACHLS8XKiNGTDlHfWnvMWGezQTrBO0EA
pWzdND4fNfy7rLQyEL0fTF+yieawp98XQEyoPnFJFQwgOEwb1z1Fxb+s1KHjm/tHjwRi/7qf/9qL
br+3hLfkFujO9iVhKZ2vR2urlXPZor7yg4Y6f7bm73hiH0Y4fRm70i6cbp9a7r8cb1dPs5wGVrRZ
1A3Q5REa85lVPJMISfwnzQZ7canUjBk1mSq77X2+6Ger29S/EbbcPp2TqqU3Vw/tEhJu+KzhDKs1
gEUvQ8kAETCJopAHZyBBjQGwTLq/1HP84czOWVrtrbnj6MfeekgNt6ZF4ygY+H+OkmFxamqDtLRf
WN3b9ssOBcqfMF+k3skFCfqq8dsai7XUFSBLDh0SWoLSdi0+3qRw8s/9oiSbc1Jun8X1npx/H91x
jrf/6PZbf0SJyiQAZjSSDpgpUHCVoXimi6bU54sLSad3lHDz87gfP2KmnFWpGG3asoe4p5jvW0Zi
xzDgBxBtxrONR9f8CysxJXyQTvG9BvNC2/X7R7ewZqCqoE7UTFdJYNIxLnxKJVEBMntbpYMjzfW9
WNSWhzVZIFygeK+FqlwsYYv3FrUyb4aOkObZ7tlruKE9MIcF+zf1PHenG/d1BNVaHXfvuqouzFgO
XkyOly254SrkPDE/chhoa+xUUkuzjucXYtDzu8Mm7fu6J1Sx5JILSYZEREQfPkcjK8luciKZ5DD9
DdqozXfGmFKbydutStppRomA6bdUV5wOtkrX568AVNiqOil+AaYokZlDKtv/BdQTC0r00cLFguiJ
XirsXowoYROmG4vz7XJojTYUnQRsue36ypaKCaAtRkqCzq/e4CaTLGrQQu/HnGGqKh/I5VNzx7mF
oPu4ZZRDgdZqvV21yX8fipKIjfLedsBTrWORAuBr7PGW7IhnWrWQfN0ewBm6TmPH3DekJ2PvNLCY
DCTqQ0NSakLvk9r9N0GUhHpYXMHJ+6mop+nkO45E5W5SZwA8oaKePAIJAtKhIvrmKt5WygmPkpOD
nDR0waeBeWzGzM/HOfnmXzwvmT6PhGi6tYxW+iogu/7krAtw7M6LvZ8n+Dx5EW0GDNVa6jD27SWP
lEuX8QWw+dc7N2DWrwoFl71Coa+yTW58nzGkt6CxUhXipaWm6otDJCtn0dyvRxrDSe2dV6W+edZw
R50b6KThGDzqiuI7beU3JBkHaXlT2bwkyjvx8D8TzILygP+IFZLYr3mENEUNQi0AYyVrDN32kZsJ
hikcB+yT4tmHfhDlis1TpnvEGSSyjAXxpc6QAwYMZ/kTdYDFyFVmBm7IwtEBUJsyypSekYlzRkOp
mROYPw7KHOAuS/iOkVhUStwVCpb30lqKtX3bykmjRAsouNMK+WlM6kAOn6CuodNzbRnmFbTX2+Dh
GyXqwINvsGfT3HHbMXCLUp9pDI9gTkCLMB0cAlGxCoVHgSG7u626XWSwf6Lm3Ozldzc7xqYbmIVP
xSt8ejDrJymJOhAJe2Q3ppTqTfFYomZPdpVwVXBu08M+sqPwqfcgnSZNS5KSLHySv7l3fYZkSO+2
lMNGP/RhSQI8WVcFWijnYgVULH7WFPMc3uvuqy3UDimocci3brMPKklnDDibb/IV1jpE1NWjhpXt
9dtPrRQ/xy75DMevNveNv7ajIChi8u1q6nh2bEE1L0uBxv6qmvDCfMB1TJuQrldDcsA8RULsqYMi
Ct1k1TiFh2HL5p3JpSIXSoig/bOa649nioKXlserk3GSrDAOWY78I6NDfZJlLIrT8vmEJQ+D7XER
ID3Bzs4oOmoija8Gg5F2h0/ApH7ssdGMrlJi6u2rMHd4pRR9VwfhZGB/wotS91B0k6kgd+A9OfHq
xT0ePk929iw6UwJ8CmWwbJWsDMAslo5RUOkEmkL40n312Qx+Rfci1NhRf/cAhssQfRTvt5XfMKKE
FUkDkRAffh7fA/wGXlmW4xDo8CpPMkkhbmpioOszOLT2uQm9TM8UEapncv5WkxJi/vevdbFqbltw
qYG9i5NFfq8j28Bk+8aypGFy02SN//BhpIaiG1/dzDYCLNhsw4Dk0lWh5+iM7mT7DKCPL76Knu4K
2jgAeJFbDQfg9HBda7SabZ8Sn62b08QX5TiREVuADZS4EzSoF8pERq36I3QF521N6Ao9bI+19I6j
EdoPdXxn53wPaOEqUddPYaPhgvdZ2YD45w0bqKwSO4L3Ha2vzyfZ3P8mONfY0jWp6r2iIxE+lgJQ
sgjNjMqYVvL4GX6Hr+tGrTG/+y0v7hy7QfpjdwNeBkwfZQAcBhTNSypetxZh/ZXfoazKKu9myezA
OakFtuuKFRPEs0OjqoK8YG0rlerDEj9fcxedv27kjdZNwrKgcIpQPy2yx9Kq9+KRKXs5rquQ7k6r
/5zdE0ijXCyFqDhdMgkl6ASluAIYFPU/iW2CxWx7C3ztmU4+dkwDpEEWC7QIpW+slFFPaHagsnok
nWQ0YX1u4xKpVMp6Ew5Fn1+/IATIAgUr8r8OwCueR56+/IX+069gr6ECQa/SCP39OlFP6pejR38N
i28ISlXK1omlipSjayP7/e5fa4op7vSacCOH0xqdJuE8/W5bBUFNgmekmM2X5MLxk7AXkgyLSUDL
jYU+eSgTZdhHH4Q459ohpYSyMAWpZcsi/K7cr8AbrDUaRW3YyxWvZciznHlgFQvpMFmLCxM27y1w
Ro7zDKgCwjjssjUtzjjbegZ8ch1tQDrj9oh7Ay8EjUocSfP8rW2GOselYGr1Wbhxh77NKUJins1M
J0iBxT4PQcNnNq43A9YjOOovzABVpkxdNIAZAHfoeNbbjsCh14ok5uDesG6y+JrKDpf5TL9mfXcG
keA223l8oOtUQpfiuAmMEzHMaB9DL6oIuO7X8jWKbluT0Ok4tiIBL4h+MNb+IoS7QGJ2gpk7zo88
qpf7DlEJlRfpPX/LmOauR1d8mMoHb1i+PEZuu2KUATt1Q7VtTL9H0MF/THe/NwGlfg/Xdt7BNdI1
46F2+4Ku+bonoSoNh1vXbWUSAoE+amDWZzQIATbLGEms0qhLkciPqdESbGJcqtrL25MTt2OQYAFM
FiOH94hFlKMBYD9sU0IksBmat35czt2Kin5s3eO/gnGJJCRkcJdzWRjnrRSOPyO5tl+thmDrkBLo
1X/HLbCVWI5w2xyBZ4y+AAUs1AOttOoEtnLB7iMo29f4nh0bm2XHuq1FWQXEpawI5ie/02DGSbsx
rL6C3x3FDrqrcZdSGiYqRpqieNLU9ArL/MeJU/YcbaeuHu02ob/lc/1JkyvIa279PkuYf4xcfRXR
xV109U/u2miOdDjcBMy+vEqgzxKgdQcq68WrDR2im28WW37YX+O2boTqKpBDCWtwr/SDuaMFMwWJ
du4Q1mYZ15CxiP1TVPIacmwZ3OHdO3yjJAqQdKCo9oGd5craxy9xi8QVIiC54YWl8IMZOjprbRib
sSUFWirt49lAhmxfPtlGX2xIZ7oPPk0MmvQx8pj/xTlaSodCDOallmoqeuZLGGZ/vebb2nPziyls
f2soAnYX20YojxxQShDfivTMzObSq/aLPZitJWzTlYe2YOwWECCES2rCEe+x+PHixixIxl9YeaWr
OBy/5WbjC2Y6nFKTJhOM7VBkeSRamnf/V0lQ1adT9xGJJaMBrvegSgZRIVSuvd26UPyQBiWp88ON
qQnQZkmGH69u4iRYzHK0pnH8cwnCSnW8BNBonC7Se1+hF+vgrrmrP0BqDO5rmhY7czanY+2isvv7
cwg5qMqcspzVGQWzfb1ycgJCOwkh9Vet+Y6MGujkxi6mBiVohCXsLzr3So2p97ONnlz93Qwumifu
Nd8Wdmjeg8VKmieo3WZiW/NsiGO7OhxkWAVvmY+6aiKvMpK7OyD/Ulew9KVTDVXs3gVL/pBx/ta9
UEPIg2Lwu++WkctPbd+K3Mof5QYUsdB2N0AuQpcWzqVWkYtAg/0RhfShdLpMUddlkwEMYnkMaeYB
eYPFCFlZAZjhvl9XQKUajfKo9nId2vghZnTl3C9z7aQqylhw2U3RUOax1akZEQKvBsE2efhNcfiZ
3E9B58U0K5VMJe9K1VLi/LzQE4edTG9Gfx3oAWVi//J13rcS6Ywlkp8GPOWBEu/pQ2ArtI4rouWV
vh9mjf8B4WT8O9kHxuxcsbmXS0hTSmiZupHbYRUe+iHfdXALe/OJVtNQJEv+IkKpE3qmnP8xFthn
VEg8DI0Kx7m1tfwyKWS5TNGjWynAKfQj7CdTgGQxvOLe1wQ58nNY+eRyNWPiYzyOJNLzJJzvJbGJ
+gkhJDP5NLtg/IoEHjnArHwy1WuUtWpd0mdtis4HqofHxZopNxIbAtDA8VOuJFJxdseug56NCt6H
62CsJuH5xr4W/VvA3i1Nfsn7Fx8GmYtjgbVgdwUwQr1DU6FnJ/pgfZRohBV5IsTPAtOC7bltYI0t
+MeHEXKeQpcyk4e9NWv65oPDAryjOtJiLjZ71DMEyFJlnlJI2TDKUo9XpBED3ritR/jGwABKfqik
ss4+88iLsozU3pujaSwPRpk7G8FvUntjSLu24zbYB0uJ9YDhivepxN+eD3MbgrJxPbUkPP6Yujpd
3pwEIoh52JJauvLDeNlbo5zqQl2iKskrNs1lojXdqwwljlugjzaXq6b8TkKAaE3z+c+eCP/VXFMG
IV+mZ0AInBJeZSUhgknFLTyShCjxfCmKys/aTbp9GCVGCCqU8TRMwVr+KU7AASpvYwNcTWO96oXl
2qrTLpGaMVdevnDyHSLTR24v2w7f9fvGNrYc8WTQmxadCb1I8QaauCXO+HE4cjphFPWSXnjY/0sC
Flfpilv4hFUxQkCCuP0hfypngyAfi1AKiwdtCs3xnQExUGOUOeXoxD0itsMUhT3IM9NC7t5bFeZl
M+p321Cor2wy5Kdb0ckwHxI0506dVrbt5GqV9h6DQzG+z5GztjJSh4QPn/PEc1IQVbmVnU2O72pj
/n0AIk50/ubuqr9Yg1iuNVIGAOkXH7OKjFdBN+uQ2ANOAsiJM22wOoQnM7C3tn+WA0tR7XUqQv/q
/4SX6hyXq4PZSsDUshhD69FLWv+j2NfGba/aqzy9f1zDVrt+5BTTZmtSWEDNlv8s66wNOrDgYl+i
jG4ggjgbrtOKF6XZ6R136an9m1ijMv05627h1Yh8TGpENvHoPbJPgc2DCKU9bTIEeqTRlTRZ5Jur
uul+InBq6WPp+pLqATWEPG+wzbPZ+c9Q4XG1MB3IjAJXDXD7St4fZ08yefUd8EHQVUOEHLapS6o8
zEzuZ2kmIy+ZAdyaL43lILIzYprA3+YbOhPFXEXwHcgl5BIKype4NtnJlvOg7W98+0RCjaswB+n1
2/7aEInhZ/jzJQfVdExTVU56xe3KIfdvAVNO3Rf+73aDXx/QJ89iG7Pa5f8I4ulrREDIDiTQWLKq
/Z73dp/TSovy5C9DGdZv2RgU3dUJkZxgF04iG/ed8+GGQ2EVM/EvBz8S+qJSVKq4bH5GVs8RiNvz
GfyVqoHz3SJvr98qKDeQTjUji83N9irsCJyw2I2Bf3T7sWmn/3NuaUcBu63dj3X420s+wbV0PNKd
en98zF9BmbJXGa/7RZ/wv7+E3wT+Z+77KHv9B6N+VhqGsjL1Byhi3+RvyxEaLsd1kgLfzo7/jxqn
8wEgBA8xO9bc7mVUIFjmPfKcZryhQBg+TxPHLJnOA5QnZDhQFfsc5PqNtYxW0rDCZ1l2L91DJAjg
x4KKvroTdvVDoGPxHA98yIOb+KKeBONknNRg7pMazu+FqOhMFLeCP4CBs1c/7QnvUvCwl+5VSTPp
N+2wVY89MoZeLnxgD+r/akXd3GWSdxRQrJVeuzxTx9k0lCz9ivOQWXAYTpmLd3X/lRlzZntiqcJv
CszXkWtnDOCx0RkM0Y3/FqwTECB0eg4+k3N+WKfiLYqKznBEo4/HIu2/+UTbr81Cb7bneXJVBg1c
SCyroG+KH6VrCS+RgTfNybHGTxoXnrqjw86xFelN7184wx+7XOQm0o6uBNZfx/Vl0cjnKkq6BPIQ
3Rxh/K2tbXNarMUqfmHqkfZIEULAo2/D5hjwghsND95kljsi1DLzEfhUkjFqoaG/z0xtVK77YA9V
7guQ0FxElMqWJW2mpLfaCjmikuRPmTlJsyS7WPjSc8MbdwgVWFEL2kQe5c16GuF6c0bYUPRVybA9
bLsfJXs/2uLulyhHLwLZtmafInGeh9OfKECju7+xag8jum/JW8w/YgERquDEwvZfUlB1XQBxApYP
DyalLkkhLfEZuiPKJz0RHCqYfniD3AhXARgPQBAoxczbXLyb3zxCszdHO0KAGL3A4YhyDS8h7Law
XswMOEb/6TNyFRxbQs9pphtf5sCbCdXXn7fsFWy1qTJ0ecMyD4veW1kgrx/y1dBqEI3MpWRH0KjL
jObuLBchebVr1bM9Au6mXOj4XHUGxxMG6px1/lsvtlshJ7QZ6O0WB5Tay5Wr+PknCVlKJ4VsYqYC
I2KQ3Z/Ku3+RnVgqewkoDoWp5wCxelrmsS9e4OuO95bO++BoRXAleRwc7/fBGymmUVq/++I7HK/Z
qMbgoZe49UtDUxGgZ0apMnO0qMyv65GfUYMXIrTrJIxb2oWXmXAhuoxPYlyUeZxCPlltK9zch9JK
pX/sMwsPYYutegfTlk1OiBdDEB8ueRGH9uageyl5i5ZacS+5hBNo0O7mdz/J9XjaLuUK7G5B2pWE
5pKa/yJCyS4thkJ4K32Bi1RO7C4uMcTwpuWwlSjmnWRFXhxk1+VXgBdAy5X9hFQV83d+H2OvnQpo
oqHG3+XJ3X3OwqROsshqeMgCFgPzMv+ScQLxvWdswG4GvQYMiMKr0VN5PS91jhYM1xjZRcIHU4Vv
U401I+pGcWJ4NEvbaxNfviwN68/YaqodDmInApGbGBQOKSE/a2WvM0Gp+08kB3R2TqPeCWHVDpxt
JG5AXlLVSgCcsUiVKuKXAVz90ajS4hjpe4TmrOQdgNsgm8bzCqxd5aU1jSz4XrvLkwGuA8PZI0Io
CAjgShkZwmNmELH/YYVMEouIj8ACIv4WMC1KfAgcPMOSrYJU4osMDV+LYKd0y3vxcaCIx/NMyTjD
CUBC0EUoUg4V+3ch739kRQnVm5bADjfg1CTa90NHnS45jjMf/qII7cIgbFTbdSy4+Y3ealT4SvWt
DaWPKhHkKn9GgHkywHhENfj+TMKIj96wis7YVD5puZjcB7Utd3Qxc8SGv1xTEv29sDBIJiGyS8BE
YAzjg7IQ3XHdDzUmBVyCOh5tFxuCLmJmU4wcL+VHZDCfGUCKGgYGp0gtDtjFm9CBvLhvpfQDE6Np
7xnhJ4y5sbpCg6GT/W0zcBikKTF1jNuwnPfDLINnBP13NnZ1kNYFUXMg8m7D+c/gFVi6/upccZ/r
N7PmeC/FBKxUxgpQJKY+vybeGnO3I5RBAKEvHlCmgtSQ8eDKXLgOQ9aqW7+hD478HgQ7JZFr/2ob
v8Qko1cWUHkqG/B6cFrc68XGKrDVmKrzbT0PN/k1aFImdX4cB14tlBtHDlGP+ge7g5X9Id0/imQh
QLkP0zh5qJGRslO6pGhyo1rOaPja5+JiiWe12Bi0HY93LUxhu8NJUuDN3aaildjVi5mViGd6aHPK
ulwyyo+rsYC1bnY+pkhUH7JN+VPMjcW5ProhJycPwXRL/qaqH4KClHdTWiBJUj28J4Qs9YpmuOon
VuQfKgywaOYqm0licY5qieCuAgoHjCwKWijcKVNRT/K3xiOLsXWbiq5cDjWl1NdtF087h3xVvFKQ
6GNqTJhdrNH/QKMWDoUQVulz/+jdgQb0U6e6OXoQ7Z+NS0yFlY4c//VvqPbu9Nipr0DELrf2ztE8
yvRnUwcfmBOzKQkghuIUOD+UY5SwjIllzWxJU5BoBS8Wj9lmkVTYHikyRFexmyzPfNx55pPd7xGr
WkBFJIiF8AZrOgoUXaUIpwiQVno7nQjVHBmaCQy+MS6CceHoSageMNcehzaZYiIUyYFDRoCbvHZz
LM7nJA0gZCw9NjZAACZm5y+jbrLTYuydbqxXULt0l7kM5Te/1HELw/sTacKbXThMoi/6qreApVaZ
q0G+bLxVN+ZF30mkWqb1UoHs14jyePvmI2ti9E5ZfLfCC0t+E65KEjCeLslLqMDvORNxK2WOBb4Y
6rPgDWMwbKWo+qqVlu2mA1tijjgRSYWKMSKGux2yLwI/cNldirP5aFxS9PrVXcwDzvMdshiJBOtP
+s5XW6FUyrakv0sE5bOZrae7WDl80xXywCAS9gSsqeewc3ZalKDaECdyFdNw8CkfhtvV7w1Hv2p3
mmBe0y6jXAkGAa2aU5VcpV2ohRlWRtLaxiYznxymTW3De0IL/R/8mGfYZVl5HZeA0B8JQfSHTkKp
eE58he8UER+dFU6ZmXCy7QIiQm96H8ykRRgUqog9ut6CLAo5k/N5pZZZt4W0I8G16rxXCIdPlnMi
syf5R/I7DGP0CGVkETxjb245qoKYIOmJx1HoQImakOKcrUftnn61kKeZvvDbsy4CLURD7R6Wo5Zo
3SJRkWQR2xq+cOejPIRjGRK0/AzRJ1oiEj0pSM0BHIo+CmCgb357pxIHazJlIKVeRGAW7x9nnVxE
PDpCADg8gLA+yyEuxtRGisQE6rB4CuV2Fs248/DSpF3YKnnb2nvFRIrR+2EhrEU4/3fcU7/d1rba
UbLSczxQ+8DtExIE0pni0gPeDeMiz2rBGerGXOLpxaqdCHmgqm01QRm2RlkpveME2h6BK6zuvWAZ
xMEmjSvQOva/C9scSuyLrBwX8Q35h8owz/0aEl/3e+kKLT3c6tb0NO2OAEe8icQdlEnC54YV+1AS
dwcaCPvZ5tULnH+4F7YJNiv+y3A/toW2exZKyGJFlbOIFeuZSyqzkuLieqk/jm2nwogyvNbMSRZ0
Mxyo+rQa+mme1NyeKhtJGNq4w1qVWaB2QtDCJ6Ghxbj+rtFkE7UMOew63rOc/UMzgmI8bf/TZv2s
exGsArUxiL8/K+Oz8nZ3c9fCOdZNauf31nCWAF4kP9e4mAGhgDZOlZ/WPZfWaz9GMIvFhVxkdsy4
mwJOx9cZ47Z/ipYWJMKaeA7+RyCqrpQtfXYpe/aupCDnFIPqPXm5XIO8tKFoK8dv2ixf/PEvgsS3
HDRzu4r1d0ovspu5QY8hY1CyZTbbNg0KYpoXCPOtBtKEGApHQE99Q59u7OU0v0G5xAbjDupQuJYA
NthAKgHixj5CkYwW213aW7+p+YYZFvrdjAeEjCZsRFwe8yLAjNqKZVVYZI90aQMy6slU0iRjUm1R
iBSvBfjUqnwCy1L2FRk2swG9wf9tRTCUccavnBoq8nRHU+Js6j+zMFPHZKLMezIaPJHZfCJVac+/
LpvcXKazUwDFoJ+nxhTG2+FE2iRbxko6QDLonaRzsHGay/oLV/xfbbLnCdiMZs5bW0C5WB4uW7kt
zQJqkimt5J/E53ZGyAOuNyH9ls42eZhz4dBSFHglbPf+nGUACYreLXKsndTVPZrcoL7kn5yEUDWo
uMbJBJgSJHvt5hQWp9rafDtGys085H8nD3v9kIRrDcdGkRSZfAa2f2XoYtTUQKEONKuyxqydFNdM
/kj0bTcNImwkubO6JeGBjWxxYDnmbhM+wDN844NJMpwU5zACz+ZEOm34SxBVYSCc9oZpB2usc8k0
q+XuqAXRV8gANPFm1rrOFbEr+eL/kgmKepgBdvJjDuC3AwcBNN8qx6+I+k3yMQkUz7RSeRDfppMu
7Qr1xgBIgx/aMSutcvpzdmpof3Y0XWbLBenYib2Wv22NLHs1UzL1ADkTBhqIOFM78nmDqh1tK6XD
IOxvDto+QrLsBCZ4u+AEhal78YiohQ8flanBRTFKbb3NZYnBy+exkCAijZzyseVUJWVhoO521UrW
SLHajBO+sgVDOgmjDQsN4XceHbflbpYwvI6PB5LjemaR0mtZpgnq5YP0kVdw8YHrQRYz4ZgoGOdP
tj+rcQFdqPqJezsMSlDmQTcPHXB6F0h3H9//sHu5ysVMACh7ytTSg0TjGXH3AB3jga/+K0XflFj7
ZLLZ3qVDb46rc3Pkto6CAvQT9Z3OUH+OqgZeLy6GxhAovZ5XKVUjtUUfx1SFtlBO/eJpxq0ruyWP
JXTas6wSiLHSQX8Lbh4YgfmnlNThBb5/OJI8Ik43scXJRRIYT2O9SEmrU/3T44/0+LsJsElkVYsD
3EvN+Wzzg6UEyishMft6lRTKHJ3aT56xkuONJTj5AtRGRFe510txppcPKr53jlbWWY3lcAkyxFNU
1KyZcKWVYNAgx4pD07d8hUYU3+h3MOAQbOeB67PnBgKJMa0AtwV5NH74ga416f42MLRE4eAVSyY/
1thAc3OEfoL8b4ls+j+uVFMSXvAKejM3JhM7GI+hEknE+awGrOsV+SoJZqUfVx2muP4joK/NtDCl
71U+6w7bpy3I2XBKwJx2+quzNITaCG9YMksN8G079lBCyiBbpFvxXBTRmItbplRFeLFvZaPqZEot
VMUE7qJQGRJ0MpJIB1MO8ulc+BLRkT1ZgsOlyjn2SWQxm6Jc9ieHv8tGd4nUV4Izp177AqI4mzC7
it8LkCgEOKsKzwSDOpLH149IRQd4dj7UHXDNKzSvLx8UDrdVkffBqOOVLoKfRc2GxarrJw+2g+b1
/Fxt8hmCKFOniLOROEB2BjWZFLwRJC0rhhBQDNw1vEg2opkMFevsBkPgoGhZpyLuQ3/yV1PPB6fp
K8Hmx1qFGfVGBNaS4xZ9f/2Eed6QfNPc/q9aWPCg2TINbfz/1dNsNJ3eTtdloR2pmPMc7dQQqoux
B5TM2kh+fa2DVM9tI3XRVIon3hKwMKFp9SoVIjzNPPmmTjkCHmlPD3ma5cjsAATwoSVjAAYoNu3u
1Cil5W3adR6XT0YJ6VMIE9pyx1LonOlVHGQFX+BDGn/WL/l5+5MXDnKtUbsXRYrj2lbXcVgajyVi
ua8q+eZ5WYWkzomS9jiO+lejlnw9xTHzRJk6Ie+5G8Ys0zEyJUYZ0jwS+tvmU0oEERRnDkZ2Ow5T
AbpRzy9SuYwew7Lgb5nkfZUe+JncpEAjX5aa8KjhX4KyU5p7d1EYw+Jrvvls3aJIpIbmv/x7HtRk
hTGv8DqFH8YwcaWiQPYm7IS7s2jsoOmt2p6E47MuYBB3bDfeEJR+cJdWXtCve7/Tc5Hl70QGavER
fR4S2SOjg3j+RZAJ1ZE6e8Z4vhG1n8wCkkNty3Y34URZ0+AlcFsYlQcKlu1qPnU8z15jLw1ZULYL
e3ERocm0CL7Kqz6RZImOEzq/93xZCcHQF3lvSPEutVstWvvezjX7yAP0GCHe04NHEQmz4eiJ31c5
gjwKW62WeYK25GrCGaKED5eARwmfVf/k+hdEZKSUFuB7R6mV17TwmfEZdF8fQmMKyChQyOa6zPvQ
81CGFSGYVOnhFG2L38UbieyxxwoQxQMrNXGM0PLvRR6roB+5XYkRe6af9hemluA0e8ayyBmw4iE1
PtMHsCbSI1lK9yLSN4M2Tyrdhssb/b7XaJQFGlKcM8R/u43IFL8DrNlplSCPIn03jruUV6HGjtle
x9MyP3SB6EH6G0+tBVYEgpiIwNP66ijE3+h6HCg2msxuSgWY4GMHxwR9vvHmtwtpd1nwMTafJjox
2kc2BfgYq1BLQsDkBFCi/ze6DwwMhKrWaFiWCiytP+O1LkOeTAIqmfg/Gv1aMaGnjpw/rC6XLn0a
b/cNw7qVN1ZXXxmDLNk7WEssRkzNvw9cvB/ajARplm/YMkvvZKdRNci5OhqVFWS8IWk3D6Zrp8ER
lNauzARa4CABNb6ty4RN2UglXQvTdKqCp+iyCt//oRq0jmQmuMdjmG7wWrype6oE1ibCpDVAY+x0
l/Fj57FPHq5mhuxIzEOzum/ri6gihkm/GTruZCJ9SZ8xAuN+lvcw5q7c4LvFOKEKofvPwhTIxbbv
+pGFdRgvYX4A0BBuBPaP1EbEG+9iqEuUvA6QLMol1Jsuc2uzcUlwuRJyDm1YEDHdl+9wstUwdrB2
8cIOa1WxzvBIpBVaiJ6s4if2udhraib1JVQ6B/LqiM6AfIh78W05eQ2F3+utgE14e99xLlvYdXuk
MFIEGo7i6Ycw4AhxkILuLs2uTMwHnQ00TO1LaExoxqCNZfkwsDSTP7mCR2/S5S2cfAsVrO8Lplnn
xRIbHrrquuYOrnXm+gzM3R1ih6JrGwF5TLsPaAA47nW6C+HdtzIqRBmj5lQpgWRVHl76lIX6F+FG
l8Rz2Zm9kHkqRsbc/JzY1f0hz1JsU/1sAsMOy1HRCKy7wpfvt2xZK3C3DETg6vfOMBx/LJHZy9e8
CCDmFGA8PZRqvF8F4zaaknem+xr+6QN9Owv9SM0oE5zQjfXbsTF/SgIMpax8bt1ylR0qRT7buj4e
kmDuK80LyXo2XDs2BG17fD/vydPig2Z76bS8sjpJgfdAmzZZSJhOXTCWYt5BORAd5oyz4RZQ5ljZ
WLM2d+5JL6gd9x/71P0h/0CZSoNprmr1vJGWHeaYnxXedq4ZSSq+MqAobK5RQOu/phmROZDwUtk/
JyTqCFfE/eGRenx3+rQBrlPOM/Altb408m3WgQzw3x5azhDXSQjOoj3YrZA+nwV3eGpY8cDLH7Oy
OjB3Q8yVwgn/Dghhr92ADnghljaRVxfyr1D8XXdkkYKsgBOvybOUzeRS6/okoXuMGP555kvvbK0f
rnyS3cP+cCJwjoj/Ur2xBMiC5NSyu1MRHzf/v8FfW3zQQcWnDJhuM0xeybTVxVKT4+8anSHqnIWt
ViGkJjln3K3GpIYDjSyCuls2PwQU5pL2BSrsxmUUeKJrbBGi+54rSbm/YrYD5M7Ap9OMF6sHDb1D
WXpTx7i1hoJOndeQ19jeoNN+HWarzfunpWNQYLbP0jxGm6UDkm5xosKnAOXzfn5Swt/A2xGCp9NL
KrAulZc0HRcv7AMRB9NAHq1bufr9zzj7dQirRz2LwWLCTI1+JXYckZOqnRjD3AK2Z363pJgZwOzx
f/GUdpBj9adtBjIkivw7GGo0dGjNg0455dOxnDYTfaay5y14GigCvpKr40tP1CXbPqeQLA63JbvT
bOvKfyQnMwDSoIWg0wmrIYrf034L1aTBVdjI65CphCzzcB+VU9mbGyH43giM/uus9Jx9mTMqlR03
1mYpn05vLid/hQbRduwrq8gxxeb99nq3kLRiQWNnWeizpAWffNQK1qJXLrvFgOS4kSwGAV7jevht
KViISc6mVSZTqXmhrJDtBewejaxLdcpb7GA874PX1VNVn6F1daxVXijNGjrDOH2pA70cIUm/kaM4
rOA7FJfbrtHv7BRPC1WixlqZ1WzC4gQQJjVXn1+M6oykmgtJ1/OlqhcKkuO2wkhIjkt6quo9IAaq
PyLgH6PPQq4ADiICf1VU9TsWns/L6cMK0crvXUG/SGz0RZcQRz7YCXsKojBkpQdLSm5Ksy2PvOIz
p7gaeQE6pJmWB9kad+18aov88864y0wIQUQ1cHe0whY17F5xWM2IeHRLUYgYGJkCvBA83yYzcZ74
aATGnzaxTTOcc7hBVeDP4KC7+vw9kkJ28ckXskczwD6nM9mgPS+zMT/uiodOj2No6VOwlKaGRRu4
6L71r7ywWjnqEsx+7IukgormwxApKiZmoFf9trih1kvRglzOxqlWlkP5q4td7ohaYq3oNBV+45+o
0ZUhGboIumGEHp5zRqjp5mhZCVVJ98hQQH7+cboKM4CzkmYDSJyVXp9tTyyWR8Llh8DCzSA7fJ63
5j/l9WynxcACk+vuM/BfFig2ek/vakXxydls36cHWTPWr9PSlwGjyVhpSkpAHFX2aprnbTDY0B6d
x+1Fn7SlD5DkzFCqMwi4cyOUFe/JIKv36H4ANRl2j5Y1SCmubHDhxyzGRGOvDm+ZpVsvCWB3FpMN
YEm6HxsmZbludbgsvOkLpi6Bnvykq9ndkBtKHKQN07E9KU/Q36Px5tdCVfvQqsiRD1Y3puGsm0iO
mUcN8hEVYEitzK72eTuZOsEaDP06Fq15Y10pAyMq6PNpbAmeat+gw0ihBEQ+yXcg4faduLOQgT7e
jG4WWmEelWb3738hKqjndKbET9F98Hq+OrB1R7/Le25zmTcVk3B5pvQB2S0R42EDF9r3ddz9VPNU
bgu3+kgBYCZ58VBJlflQB73MywhcA/D9wUS/IHPOSF4ab8wdps4xzQP8jwx3tA44eUdjneSErkZ4
EQ2lQ74ivZKnskIHtV6sZB+ePbTDTEyOMSBbW01/uW3OIq210n3RrSox9my+sw8gCfaeZ8buclJ3
Q7oVSVvH8ldn85rX1UzUxbkt57wt9a0mSqGP5ez+mEsu/qPaFTYmIwNtAN+XmYWG+Ofd1V36YqPd
/PdIZ++fmU2jvPbEPv52CLIwiTA0ELmCrkmnjCJqy5kV0OTgim4TcG3Z3L3A/c5WxsuCwgLCEs0t
eBoFAhU9PVhMIS5ySTygxXDX5nTJ7tJjxTu43VpmBU3ihdE+y3c65suWXJ6YiVoqTEiDGLGvtgeR
WLKFQaPWN1ewLSchZgtmFpp5n73yPkGxY3oJzAhzz1qp14XWPv05uC77iEIWJx9Lai3t3Uq0yUCX
TC/iDmGaTTOx3r8AUa86kMkPdVfRdG6eU+bAdnF/IFEDFcGOSB7lhwZ8EBLsw64/VHD4ePNavbqR
d9hotia3n8soeDKDpWq6ywweWY7ey8nEf0k9s0J2RC8KMNSQk5QgbDHhTilW6YAo3SPvwjSCPQ8e
Dds46ogiGC6lZa85YtnMjs2pa2VhcmbcTMteL7UJB5Y59rE8ukB+E4I5gxdsoiRHWCa3PGGHW4mn
cbv7/Isylf1MUktTMcDTzOZ5OZ3LEl4zU3IeoJTDpMaEeHr6gaumS2kx0hozNK4g+Q+7bdleSZwn
ROJGrX91w6nPzZuA262SN8a6X2XPANyFQW6T5ICgg79Iq/o575iNas/4bWauRRJqhq2qdX+e29Gu
DbAJGqbJosfAdM/Jn6ffxvUP93VEtUm0Vwp6/p/2swTQRlkrnEeDiy0t0pYEZzQsMj9iknk0Z036
6Y6ZJfPIvBh1nbh7jJ2MDmia4dShEL7OKH08VqWiQP0namhhrTRBhyyHOiXufi4T/zBVbQEvKiIn
zExGUfhIr2/i8+CV8RPgJShu1TfPAFb0op9kctWoGiJMCVSgdshBjddXWiJYxnrG9V1Hti3bns8c
Y5M2C8Lni4oPPK3hkEoOlJ84F2sYM1yUAvfH0kS/TdvGyIyEP1x0iwFP6NERXv4yWMiEWTAymRLg
0OXskJSsG0y2QM3jHq6dRCIkd2kTrlydaVjCBod3GQQeYKXdT4iq62lSX4By2sNEIWCxbS09cUEb
XrAmUs3mJ+slWCX0OcEK/hSYsx8klEl9IzTm/sj/Sh+Dr1tA/FJ7ooToz1sqkLP8N7mwHIIOAdIi
Bj13GVouwjjsHqco4om5ZSy6ci1YWZB29HpPDkCquU9+2DbgYzv23SJJOFTrYj7jd3TBesToeC39
RzkZhJ99zizHt1l2k3c1eIHLiWD6b3fvlKJiyxQEaYksRjQgsDyj/lF19HJgEq7jWm5fM8GjICRP
dhNV+2VT1aNG47pvAsY0lTtulT8Ug/PhE7L3+NFRLmol8N2Gmk4uq0YALcQIPyDGQeUja1oICCk4
VsXpU44kvVnM/C0xSNn2oFoC7LHp4U+7XB3hlYuMEcN1NyNE9kj3gyE9IHyilhctSGqtmIYywygN
LIt5UCSqZypGsIvLZ5b9hhmuBVWxtsxRijgbGGT/W1tJOVnJt5n8F5o55LTjCj9Y2rE9lg4u72Qh
oxfutQ3T8vjcOdmmsJAZlAtQ9ywANEekH46bArTnQPie5b4PPCbmfC4eLdR2qcnn4AGNkJBaWwXU
QmHn0wcO0OPQkLk1/NEi+PG6L9Urbhtgho+j8eLZ+kAqOqYY3NqOItIF+03twaszoyRfGqDWom/M
eIrWOeaAzd4imOJ45AF38yOaRLQ15B23Udtn5nv92tVbKyiANX8ON30io2eFeQyilmMHkK3wvem0
mRa077U8nU54DAXV8YaCBXpAzJmvR5f9P+UVBsV6RgzxmigHJcOJj2VElv4qJJhJPedJzMyZA/te
i4sZQfSmlrbOaiJqGxiIoidQSbbhZGx1pbU6sjonJTObQZD049QGfAPGWlVHASgpUyMTYMOZ5+fQ
auTYcXVZv5dOqYEtlAo2iryLY6Plvr2Jpev53BNRFuZSUBGSMJDnsy+sPCYxx4QepnIVVMfyci2r
gw4r/XDwMCPPZQrnzgy0hrOy+CGZnadnSa2vNm2yjxqCt8JYNOmf9TXSOTj0B3nQj5eMu9wRXhsE
FLLq1Npn8rCRA2eCib8/7GYGawFjuobRV0Lh+3jXPFAqFLjMh3lMzX+CAoI1luvcU0BZV3aIaE3T
/v4cQZwH3mdiapNH8EEvu2DEVGNjblbLqfKSS5aJ/Xg0IKxuU9JLwWrAOF/WkfNrK5TuE9wEwing
GmdS2XgYauLe0Ea+dnIjxehl3gPWbGbONzN5ez15xEHm8NnKK2Fsj/1XRp4sUA6BLUf5HOq4Cedr
NE5V6PMGzDTxeSXAa7+9DkYp6pdK/3uID/mVe8ZmplBZ7UmIDjaeFDFvP7HoZKW0VbfCSccdlFcK
rzRK3yN0f8ylxzGc31INhejtppv7JyNRi5iqJUnpCtZZ68/+gw4yDMHMR+9NvlKqPmyfgOfE2dtf
bFtkkdY91sNSQ60n2hmsHcMSgBSyFqAv+O6o7odbb51VjCI5sIKcboB3GlpO40c5b63HK4GnT8vH
R7uQt9lC19xKPghLwuopD7AIb/R/GK2Qf0JbreKnMb19oBouYXV/sDTEXlNitMp1J76zZpGrnQI+
iMoLJjw9NqgYg9OKoQSZ8s7BS8KklshclXhWUwUp+AsdeWGSAcd4pLVJNTAwsLQXv+jaUIcZCy6i
TsTFZtcjtO/yjYHZ7nBGXzTvz5uvS1KHOZDKtbXKBLXP4PO4IUJxa5XHjgsVbS+hIfMyu3SJSn4s
Swsv/5q2+kJoYZkIl/wsB/VNUzkrvVIqxd7DD3MQ0R40WJ95XKJ8VClztP6hYPJIYGzmCIEStQAB
Ux+5kD1pLIB9ZfGCoUNqdZfLV2JJnw8UYUjwtFs4TU9EawW2YcN8pEfAyUog90bDHmEAGeR1/l8Q
vIjVM65Qykh2UqeNjUgGC2CKveHwLzYxyna2VoQOeHYpGaVF6QNcHmStr0Qze95i417OFNbZRbPe
aJTLDVTEfmOH7k0aX6mQYUDofzMlHQjTr+V4590ltv41Z/Eo78YliM9Y6uo9syfL/fhj0La4709g
GuvvUBClqZlxcwGeFVWoBgVDo90jiUecMssstf0n89r6MkR/97KtSgwVd28DxzFB03rY7uyjm9IE
yqFu/ynU0ggpssjlJIr9SlVlff1Zb2bYSr67MgzePd5OuJbVstOTFYuFUhbOqz7aurD1Hbq1lb0O
eN3ZUUHHxrc9SEcyk0ljTqZEIp4ipEFE91iHSpihSH/Lqy5Z8AhhHKTaH9b8rzRI+6LvF48pYqB/
9SoZix9ViXrFN8BtUdDsxV1eMQoI8vqe9Nif/pkonBm7K9gF0ZELUumFLg3zgUd8Eiyb5d0NKK//
NSi8jFeUIwhf2yNTH23sKg8+vX3ETbXbuAR+i3QGb3FB7cC01Wo4NQ21CFi2K0EjTWRCMgNdvmJ5
Z+cXLnU4pWZSrqT/UoaFoVdB1B6S5lzR75fShoLC304vETCNwOy1pQhrrugWMy1SvpptbFm+aQ7J
XagsIkoApNDg1q6qeCa0sOGQFeTgeotO14sI1dRA0tinvyJlcwGVUqe0rK8vUJmCz/h6xNv4wveu
X0o+FKrUmGiJN/9tV9fg4Q4dUoSOvvtHtruR72pgencQddpmis+qZl5FRmBMvHfTuS8WxUik6pvz
btswK5Shx+sbFw7O7GB/M8YNCrQd55w/tUWjdeJZhuxEiw57dvrQ0zKosF99kzi2U8ma7uSOAd5r
7keofjAEcoWGypGUVmlSp5j77jC5nG4altLYlzN9W07gXDsaIdloaTAbvNxDhLgOMNGW0HuYuJMH
l7y/d9Kj8RExbmVTGisi+LXgfHMoQYFK9B44LpwUN5zw5U3+bzLKM0KZ8j2QTn1TdyvR5j0OKeXA
xL8Hu8BwNi/I3N5PvRScINBoArS/2qZtSfuy8c54gUNTlzoVqrX3bYBL7bMO4rU+h/gGXCfaMo6/
MHm4pXXA0JnkBT/imkNWKNS5IbXedWvWF4wd+AT+EQu2pjl5leNbnhkb1ftJcyPDkXyJ714ryNEG
lf6//EUpqmxtyu1YXEMK8n7O4L7WC/llvBUoKPSmy5+5tetJYD+iyQYwIO2WIvpCVVpkb1TBYE3D
YbZmYUAOrb1hcPMkAF4P4O4IRUzNpvyDaPyB+nN8AvZqBbrWgx5PXI5JN06ELAcjAPN97qhXhDHB
TUeKoibWD9Ut6uoDMLm8B9O7WM9K1LmJ3FQd3DNrlFPZWxyOXqsbygGussjDg07xPfxAvucwXpQd
eoGkvFYrbczdC1F5W9b1GwXq1oAw36A7RrM/ancICsgZkD0DlsUw3cic/gEZUC8EIPkWfH0+Ypdr
mExmoy1osMEkD3Yg7urqxcvIo4NaIMb9Tdi+KRSsUbrux6g1OqwfhBmG0SmIaJiFu3Q6ccAaSpyS
XOrA2hBdTSwU0nLFbgfnHzugl7qRFLnrRy9RBBlN9BrnPNN5j533tHRast9GhopwQ9YwkS+TwjFQ
gFYiQYI2qR3D6MyXdsMZO+i8E7SyYrNo2AJZtcDLkXRI4MQVaAtXU44+ucQi+W/+Ny6IgWl3IGDu
a+cJ6FXYpA3wFfYV7vyGBD4wiH1dncFKgXkaQW/SOqiYeurs9rMqep5myV9Xg+lQN5vX2Ab6zEFk
pWH2oZKtgbl4YgqH5Ec920V1gqNxhNh9qV+LQPEX39p+aNRpYiurke7APUJxpAuik4si3OdCACyo
rsSrZ24iT13H8H6QptY7uOk7t5ttex5NmmjIgc3dC4yAyQnCitj4n6Y0X6HrTJbOKwJblmGiiI5a
afz05KKMlkxreXBFOn9SwNkscGCFSQ1L7QMswBs94IivI3Bb0dZlg7lcC8f1//v+jV5ylKMEucRu
5DlzvBbabBnw44DGCuDiIu7ATeiWxXgez3LzL7uQ7Ez48ca1dtkfLtZmUoR0bW9k/VhoJYmvTrrT
h1wm9MBHXun2LMxwijVe7BAT1XZ6NV63rjQKJfjDsuceDGBAj1Q/9um4gWnjP7LTTQKZeBgYA+uy
ZmkDunnwiAImaYL5x/rPXkFjzn4KdbD63WUF3SsXtpXbgnz4/crr3JrJM+/xhQ7VIyPUUNvUbCyl
p0pI7mTqGxWjR5StFJaMwpY6bnAm8j49yR/QPCMhbQ3x1NeIgLB+MdIAFPblBZ5aPn4SlVH54PLE
/46RGy69omvu+U9U515ErWigSXXT9lkxLCOhxaowo1kJwQAPPrzFwuNzWVsKsS72o7z5RUQmlD9Z
/5vSD0uXYKN2NJViL2pb5Eo7a5poLGjrhFj/JDneWVOYm6JP86x0cxL0KFXHOhXKG5+jo5Ny3/Qi
lwvh/DlP7VrcCuUTRqSFNspNCaVwhp3Cow0ED99qFN1Y8rczEowZq8wHtx7zwkHQvbUiQYR6qDgT
9duP5fmAqkoyhHau+bEHnBFlzzLau65uFCiXhINznIgumkZa3bV+QGGFRggtwcnds4QJadIdFub8
Wj+Orpk8zHz/eAEcVMUUZpDt6+V1LyVl6OoyXYH/gGF4zIFUorr1BLRWz78Uecxw2BNaG1YPdviN
8Et2CCkPpetxnzTrTrYZYs/kNdotz7Ak8/e6nMyNv36t3x6MqoVjtm/itYM6L/X+QM/bBBrtz8Sq
aU/M4645iBK5JefjDOEFIX//i7jHPUoGAWc1MLjhp1RihKaJ31fvQrgiyRheD3tPY+CHHYRkn/z6
ufigj57swmO7essietFG6CSUpJvo0mzpygXFlC2noiMesnv9gKGZqKvcpoJRShURzL6twGavVdFS
h8Mk+s69tmxl9I6O3Q2Q5jPQjIoVNl3ff7SurL+gPjj3J3BYr44N1erWSGI6Ohf+v+V+gseoeT31
zetR/o6GuKK/OkWNgy7j7uyXjVNBP8iB7vJrwZ+Y2YmeWjunTKMoriyPZblYWnXwlTUcL1Ofs+vr
4itD7VgtwuUocWWC54t339WqJqN7MT6sIX6Ehmoi7f1rLkdlhfoDlNfjKwxi3gRb1eVuVO+Wucxq
BRPyO7XlFxX4kVrV/hrc5l/Ot27Ws+y7lypkVax58vzkBhJiwMyh4xo3qeKgsKcQAXdgyCsVIck7
wPg8O3fGYo8e1zOl3X6gDf3QE5vA63fWr/A9PBhPqxG1Wn4UyDtzy7FaWDFHfVpi3IAT6K+aGVRM
huj6JD7xxHMlLy6o3zpRlNLbGuIKMtt2psnhUgh/KPJgWeL8paF5gkxCBAd/pIPGXLc0UbJJOp/G
YjPWMSsMfW1lc2edXf51+0o11+2ttnHX/PLXGEbHvLIK4Dm5aLWow/0UWt6mtlQ0jGSgWqBBtki1
0ApG9hSusaR67g7qDv2FTfg66YyKeaOt5tXkW1T6yxYZcaXtgfxDY9c388nKDFANNGMFQzAZultD
/7pdufoxsDeJ+Irk2VbXfHi60QF+JuSp3smdTEfK32lMrsu/0auWhd0kCPZEteGC5UvbzITn05jg
mD+SiP2dqdykUOxTlVyoEo5Lp55xNb8eezhPaZf0gI6lGYwgWi3JlXKT3/NjUIwZjSXY/LpQJLqW
fxdY3zY7jP79umVZkJyss/ZygoRB/+H7KosmjFGUrgPcI0lPR91I3dXtVxfinFxKvujn7x9wpc3x
aYjpu4zWdEier4CKMZkZDVEtGIQbq+NxRc4LGOmr0eA7AMOQgBf0uAcaUD5QPTv4Bc+jANMLsIZA
gwC8tNRm5uSnnVSwcndg1pQQE8/o7QaymfJa5YBNwZUA0v7AipbqFbeJHJl1pN+rlaAtVJ4f/igC
xUNTfbxja80sGjL4yWcGerTiMG1OATnbypumAALhRCh2v6nM1tC0oCc0r8nc5lxLYhBAMR08Uu5U
lylpDPA6ogTBhqtqprvhbqcGW6zL+dOJzeuhcVRZbXWCw+/5EcexH5RG9Zq0nQ+XiX3OaOZB/HJ8
duZA9swDGvjDlbS6HFV504plgDLe5vos3X+eAFJEISoYhN4pdm6R+UmNVL3dajt0j+2x4Fe7ivF/
La960WNNd4p2K3mRfmB5318Qy+vfxk4Te/DnNcYwguf7nDWGOZkVB6tdoovGPiEUsUc0F0ALWP4C
dUhj80GkivouuIOoJPdZZXzC/NdM8Xde2GybxflSdJJeMyxIhmO76tdQ5LlOUxWYDmGk2+C57Tsf
J4oBUv9UsCxT4yl1dC7jpMx370EAoLRV+C9gADc0JTPE8dSuQX1FpLpJxDd/pL0GcTS1/TNhJiTf
gUtKHiDapTL0IOyEt1BNlRYeZC9fpvV41sBNevupZC75Li043wZ1m8jQ6YwLVq72Z3Vrh9DayGv/
LzWAJO7HrprK3VW8o3aIIWBvXrAb9ztF5yLafvDp82osLEyMNQx1/FD/oXM//GUOhfwWWVPYj/2N
q8DrxhTw3AwNjwnuCVA0uBfjzGzAVg8kwUHYitjyQEYRs92rsrp6/IeNog1Q42N7Jpt8tsiFA/dj
bAKSWqwIH31K45sS7gdAv1lDZXaigy+Cmbf/t4/waV6y9Fw87Lzz3OOUnwCMXRz/JfcuZvgmm3SM
lqGUs39uKoOtKSG9D0FC/Swu59zSQqiTwQyG4BFaT8WXNjMp/KvODD5D5MwrYUxPLedBq8m2oMDF
f2YyGFoUGDj3HQ30NNVjAHi/V979AuU+DNHjUHpwqPuj6D8SH2k+oj18Vup3wldsSi77/+RJOPvv
hcav0gX2X3DQaD5310TmhcFJkh9o4KKUo10hXhVA83gcKaYzQHT5xgq6k6ekUWv614eP5WAY1LyH
MUra+1l1QpVpxXaCzrhBIEBA71BgmWYUu4VUgzR4jZlcT9qNtI2BLVwdln7VCA/XDdSZion2Uguu
dofznfMF5OGF54MBi1g9AjowhQ1thzdsoHPdjcdw1qSJeF9IuHDOZAHvoCOZdzW76qN4CdHX/iCh
7b/R1zseUseiEpvyn6d/8cXyu46df8dDQAlBi+VrmPGhA6fIP2JuU+Eez873xPGRkvrm9yv2s1CH
Dlh4tUdSoTk0mu9qpPOwpSy1Xy1J7GVVaTRpyfrPM+6YI5R6NWsbmJB9BvEOCrjF+6ovyT3hyVJU
OsobvYxiohZ5pAO/HqwsSmT+Nbc6/1zhKZ2q8KSI5At03KOqS5bUlgA4Jfz0zmLUhWrEq3dDGtip
8pvnyF45wN9rmxnB6Q1jtqfAWBTX5BMXT6PpJyu+FvVa9jZprQa8uMQy2gJokJyTBfTbU28FK8dC
XUsQiSkXWvcjN46JnJBx3rvK2zuzs+RZpd0o/F1xpHJn6SqbHqJf5QWlSg7/WupeT0Dj9OdE8ctv
n4+cqYh3Fi6KHeCGZRHBbk9Ym8wsTb554OPZhSlBrOGhm7Ny9GFzFbBsVW9FQhaQbqBIBV8rUZ8g
EEenGn4a4I/SnVk0y9FPAiNAuG8ShLgtW761LoB4N519O69jJTgBE+0koXnw4MDnkzH8D8krQ/aL
JTX7bJj6blxnb7vxZuTK8RGLyXM9lQ+Xh/sIs6jAVqFWg9F9c6LbNxWtTdGyhTSEDLBsOckdIddN
hv8jJjndcumH2NZ11+lqd9jkd8URf4yL8Cq/9q+gVyA7I/kRZwOnruxKefgsxiHRua3KG9fHKfRo
9RcSwrmCxaaakctHxZbF+ZJU/ocB/XefX/IP7ZrN8AWYoPVHpp0IGm17lsiN5nXVl47goFe677Ag
3Im2rpGf6h0XVO1csX+C3v0tJ2q6fsXqEp7Pw1aMDgwlgaEVaPYeSykfkDv50GMUWfNwar4wicV0
E6k9yQG1rHZjwa7PYBrxgfwUBiLPVDEc/NRTLGG8OY7JZeD6E/15ylRXW1lzHmq2P1yck37faFEB
/XQGxaTF9EHGAdUKqKZitQzDUGalucPhVqTIJ71HOw43O28S+2KVQbBs3arTnwVeabnffsj5iIea
H/G49oAXb819SqkFQyJqrAYxccD0BVqS3RZKcSu6+648yV0wj8vwPI4SKWMeJI1jBlTn3oEDAv0P
6iUOR83ySKEmdOmmOr1eXLeLClA3s63BBqQ1ULgHo7H4pgRGfM9X7phmfXg3lW8Sic2AQn/pZUOS
G4M8UCQfawPjD5S2qfxi+DFpx7U0Bq8LlsuYDyH+G2CG65gJyngBoEJhGHBbNXB7H7SuDUmi74BB
wqZf+TOA+G/tKcMA16wMSjNgPHZzMuczW0QBhw1Bs8dXMe2t0MpVVb/V+0mLz8FuekF5prM8D/zG
axXlmkONZ7UU/7Zkab9JAg72Op1Gs0V3SbuhLgg2hV0+6LjB9u2XmUXWR+018M7BZ7Yl3d2owvqg
OonQjpiBzqSM/I+T+WwgZnyEDijFVEl9v4J67X0p6SLjsYPKLI7bGnqpfba76HTRk7mB5DrwgZxo
sWhCd5FRHFJfnpnRAMj88WPMj9F9UoGF6y6Y/yJvwcnD8klcjF4DwzyB7PoXn7tr2KgyUYZHdHpf
rIftIuvHgDke9uNk2ecRoXdmzSvITUAPNwSSYsb9Z0slPd3zLhLvQ8QchFwgai6KhKzDZAGrH5eA
uxd3VMTZOHjWTpiZ/JL18PZLI5Wc9sweSn5D3lvHXQU8tqKxYtdM3YqifJcxB4ovls9O/NO6tnFe
7TM2cl6sGhO76Q7ryZiyCkkMxC9ipQdStKT5Di8aDoGj+ukdtihhQDhPy+nrDa9QZzZ4SuWadVL+
FzSeJxRHUgrkHU/5pu9x4coCwt3vl1FhooCU+wEJuMbuFiaM7RGzOgHyyR7Vid4ZoqaQcmOr0EL0
6ZejpoF5jelR+zmyDoP/y62DaoI1xP30ql/iVbU2JZjLXyFE1/bqG3sHGBQ0b3CMXbEeLkFfsCyK
PhCmnzP9cK9cGcQHwogsKESeu7OywkgibG4TSomEav+0sbZcoUEjQ43k8PLZ1FLi/nSMG2ZLPL0P
p2J8vDpuoGTopZtXszAZTGX9GDQwEoXTAv2iN9pHk24PC3i2vsSrjelnnyjU2/M0j/NMDf+C/Yqu
hux41wXtttOy8qc71SSy0qjqwiMfyO0bfTU6Bhbxsi1wbpmrLm9l2pbyGCImmWsVsZh9qfo0kWG8
/7SnAbNnxWKPSxjUBB6r7B0i5cMtsiXntpcJFAbE8tY/SOtD+x9J1a+O0BpO/IOTFZJE8f15JOMF
lANhkFwWl9FHSRQ+z7SIz6G25ZOqDHGSvDZ5tsSwFg5c6snpUenF6Bm1b7XruEQ+fBEu7kKxEM6f
7kNvuSFmslesGT8jMCy4G2dhjtrc/gKdW2+yo4DGs0TQZG9eufEMzVJ/0joVQOUri3K+YsIDq4y2
g7KV7fklDvIo2fnc+MVvNBV3RsH0bPaRUrzcuOUyqnsGaSpx6lboTZt3Kbnn0n1WybQFjTZNT4wU
tyTmifywHA/nNM4TfPdfBoOorD0XAxicYB/m2s2ZaMGP9f4plkxTn2OSd4XVoK/0n505tpyW6hbV
BgL4zJjhq793L0NaNpcZgFuRnxvxzH9kFLaGTQyYaJId2X7NtA0Hxr4VcDAkovfQ16cr6O/87kra
KByiv1esTnnGUCg2AAXO+AflIi8oce6Tqt1TNz48y2GEf8kUvVHWBDDbiRH/yNnBNEakujdQ+bB9
+m7+2BU/QtmUOSFJC5te0AqtVXzxJwRaYYgdO6P5BAdaVb/k4x0UJNpJwUIk8sQihtOyLgP1XE2C
XHAvtGXj5Wt9piq4XE4XBVLQCsO3wd7GOzGMhTlaeYD+n7tUrcnuEs+s1pQDSA4EtiyTEwVV14YE
XH7B91R8z4omeFnB6STQorUhC9LT6ehxynvbsJBDXlB240/bq136S+56wT3BcBZ+qTw9rsXGtBN8
FEdLD8cpfIeAeQNHbUKT3/DxWIq76CFiqMm81TRe+WKHeFXJM+nHYr1pqixBeT8G83JuNSfYyXki
EyBe7GDoWXroUIkEve9HP/R/ojfPZ/LyVGGXoDem3yrEABKiKjTfza8u5rjKcUZpDRv6UoRPQJCj
trqQi9zpWB2ATObwSyW9oMcSBUKkDtit2U7zg1x82WBHe2Jfvr4IHjmgwDH7vPn4tw4+GC/R4bBC
0I9fLU8zMmA0ibKhkrVMBqpqaf85/oOnjbXJ4gjR4x7StKb2FlqlDUO+Phh+QUz0i4oQPrMhosaO
7Hcm6Su6WY7WwzFe6+LA2wTEdkwYQl7YPovhIE4mbKDk+sbS43pUYdF8Ty8FOehHoMHxpVFQ5EGo
Q+r6Er5AtAUw5stQx2tHcKmSPi5w1MpNW3AH4a4eoorQGkuSPvW8eaO3/MiaI3r4ZqKZKoEmwxRD
lDA6GfzBkCbw2xcvzBSsFiS7bhXCMwU6GaDwZR7q+ZorIjP4f8FozZjJdsgixGnPLVGXFgXJOT17
SQLgSjZlyi6G5AXSg3q1dO1K4roY9JPzLUmMZqDdVkX6y5d+ML3lM28RpFTM2JvUukvIfuNhoxS4
v2WiNwv9mqAhLb/p0uvuQbEIX285tnN91Jl2DMaKuHnl7dWJPJVs2GbHNwpcq6K1WEUIGDMyV2yD
oauY6owqqEeTAeGYYheYvF/lJFD1djv4Pzeo1oc4/TQjyLnDN9R0t4XRtnGqn58H39y67+sBm19q
6IPCEnDwQ60S31PgR4XnNlwuM6naSQUFqqZxyZFMNDeJOmQBaRqjsqiW1ZkPag1lfY3yv1xVqDoo
Tno6jsqGlfI82exP0zqiShU+d0TH4Ucm6QkyVQIxgX7tkYFito0pB8O5WxFuNrUH7aon7EofOHo9
mAs+zSixaXBuy166AbKrfhvmQgWKzJUZwOAPInhXsQn3/tzDX4ccdKL0CHXXmt1oqdHLFZfttCh5
LjNvWT3wVlGyL+5zA4lz8YS7wojrzSk7fY6rGN/YcN/jaJd6LTrxVSF/y6xovAvlkwvz0BLREjjU
omViSJltoq0OL7SB0YhSTR98lokLCUzPgIVgSS13akauWAvDg0HjHUldrGZfqATZI+uTNjNEhAr9
8GoEteZctGSfdJ1KNYf3RIth0RAQDFBuqizMgdCQqzNYXJ7tgkbnQsVipnRId2eWVEjkRTIXyzFm
d8ygeg37hqIqg14Hh/u0xIagcSekiG/iV3E595WEYRREze3xHvSRY45yCznDD+f0OC6dpKobvuY+
iI/ODhSyQeyXHCrLW98Qvh5q+TrUQ8Oc6FHlu7kqmG1M4UL+6OhVQ0LNhixO2HEbq/W0LU+1VcdM
GF5s9nzbOLnEc8Vf/WAv7+bl3voVJ2SVTFGgrLjhKxS9MTMvuvlVIVA5kj3U3JdkQCNCn74MZweJ
h3YRcY8AlhTbLaaZgOtbRtC0KQjqWWbM2xKNAMYVNpG3Fz9EfAaOkWmK7JC2jmzk6aL5a3lnjJl+
bR2295Mdz2OgcLB5l1T93n/YbccjKCqRVM7CeD/mNCLiRIgXSI0BvTk+qLIJ8umgh24CsTnfLOrO
hl0+ZoJxYB1DXVPznlfBRcZhk1jGtV0zipc0Mxf0V89+VukuOPwVnZpHiNDbsJpGIXsrpSD9T4H5
rMi9D7VSF3izTs38J1m9vDEoeCclAavLWAL+G/Opy0JJqS2Gv8j0Z58a3LBgKEH+UnXLctxyBPZO
gZMIOjsKueXuZeqc1fIg++czTriu+++bvGeMPoIw24h2nMmPIGkqHG9LsbgauFEiCbYWlVXRMt0B
Mt7r4TdCoLyHCMQDN31UYXJGu/u8/OZ0IxryMOTi65bquvSDcDA3FRglUsRGJppCZElpDsLO8lw4
CJNVwt6u00SMcr9pJRtyFtnMhg8xvkFSduykTb98EgDLU8s/ldojloVAX50JV6nO87wmHYU44v8Z
vQYmbmtdzBhsDnODPIxHD6hQNeWFljBO0cHTRK1L5qUbcxEGpLTFC5fVh1BzaEnhi9LdF7oHHuRr
RBmVyZ33AWoWrNkk7GYeOHmMhACQpEHWdV/LvajlZPXWT4B+Lbl4QE3dMjnwsLsqsI+q9VrIoL5H
d8FOTD/4jjfwNXBe0dTXmZvZDmAl8/s/+M1d3zhJpJG/jHuAfw8cPAmZ48fGgoA55+m0qPEO0d/x
DzefRmhUvjJvHxShAeGpSkTN60+D6tT0vcR5PdsiP1JUNHCA/5No7YHeLcKSkhtbNM9M/DiJFvaJ
rJkQgJVRqlhotuM6U3JEbGslySTTsz9T3/4tXafx4Gxptqh7kvOjPtINVu6KQYw3n8ezuonA+PPm
32TNYG41Mu8SuJm1/cdG7xWhgA0iegysMiONTYOPEcZAfRk759EzeYOn4TInlC9R0gZkdDUbTISJ
IZ2YZaRAADhQJkUEIGSp41ySfKOKAo9yOaK6XVe4Vmnt4IITc0AGDmmF+vBJvEWxrhO/Qm3ProEG
/i5ls401eUNV/rvBfBp+3+JfLRBsHW0KUC8lkGmHHgKo3yTecJ7lMWcaObTKiaOlZXexp7FRf+74
dClKyJWi4IwDS51E3l5I36tXD+LNrw21DLBJ/VAQTG1jJsId6qyDSp/zWsS8jhXBvOMALF56PlTo
sam+R0FLRmaUBXUrbgzfelJtOIFK4ca6yb5NnoPjNGD7nWOWaCRXEkMbT4fe7W6Cy57a+6IPEvXV
WmtISkHp+lH6dmsnqoeB/v1g+o6FJFd/Ol1UqIg89Ae/L5FyKyehy8ZP1zJigepSuMose1ERUGtz
y0AFJ1Bn9XOXfAmUOUB57ul1RYb7UPbCOCLpqgpxFord1Ix3rrCnUjCySL7E4ddvAMLkKZHotZzA
Tpl/KWKRUKJbJTU6SpHSUwDoiTkNX5k+BuQjEBIcYWk5spjWlMENGKuCzSMuSEhxE6aXsYb8ohhM
8lKlU1euutACi2n2sEwrq/UNFZ43f/rAouoQVNt6IXtbbRKOhCpRhHvvZTkIZpBI/2fOWqFq1VBL
sV4GKznvvxNqBa7fQ/EP6BRr2AFMeE5P0hvSFBDtr6AwjWBHN/VGvu/ZympHGp9Q+xIyOsvtuvp0
CHE+A9KlfjmwHheJOLhbMHzKD5pxpe9rQ5JpHyFPTZqPwgvxw6Fa666L7l7Dh6hQP4Og6S1MCA8T
aHA6LHaEDOMVMeADfd+29EqX9SIRF6Ds8sbha4hDKejGh5lsBi5pp2GJugoGZqiqLTulvesAx1WZ
ZBMnp1JFfIOETWAzhvLe/b5cu0KVKAfQlQp6H5Y1/XAAbGAgyTXm76fwIeRtEHQgUmQ2XdK9apg9
tVL1SPrDXV3Ahjmha9FOA5qplysEhgv7BnPtXY4ALQYYaH8DYEJ/E6z1itOPqBg+N56oHxku7m2U
+bx4onMUagVlz5ZfxrYfPHyIracJscYDxwaSJ0rBXpqnkgWb2Zc7vL3D/W34ZByjY6sazTriIJbr
0lcemkVnc+9CCUQSIqoVdQ4pvzU2LXEelelcUP9kYggp3Bu9v9JcGb32T1EFjqQ3nr17w1Ijde6/
U8UNGSNX7yLBawW3zxQHq1yhKOd4gNmRu5eulEQNV51kfDVhLgjm+N6ly0SIRIOYssxKRK1b0488
VqyEYCXlSEgeu/1ARJo0zgrG0URRapJ+BLTGdTUssRJIEMjbXndliZaKgrL0o2SAPvbmmw0ucFva
Nq5VaMnc1ta5mAnWfzwtsIYpxFjDUFwmaituMkC0Q2zc+NEKsWrZ8w2ZpUrrKUszyZbuGaAMRMIu
FxgjCsbOHQhFR9Plw/IU7WOWRL37gBZt+NsolohDHlGTjzLhrcc+8VGdXH7JzvmVg+eVXEKIxmDe
aP3Ew34bys6phvdUpXhlO+WtIcRj2oOzA09YzHv8XwHGiT5fVrOe+GGhGiRtatrSYaKMW8VNXbVZ
4PMUPUSLYz668wHpCe96CtJ8BXZ2PKVCGU6HFSaFb/s18bqUDgjE1nLUApZ0+eDI65JJ40IazaGe
mgo6uLifZ/wWMlAlZ0+h3PiIz+mgohyC1MlmyfXHRGRw1+oBB4q+LhQySiUc1wxhvm8Yz5BJV9fX
wZQcpJpaU+uRkKUET/B6dG/ovdYWH6cQIP8ZaffQZiZHcILPrdDIwQuLMnW88Dd9HQdpaNuNspDe
1GDLMp6/O/Zk/M2c4HHC9t7gjyIILQHv0jhYypcHrOZXO6lJiFMse0DLlTJwEAc9XsxLSvbkbVn5
Eux3ia4i+/tBupwt/NlnFeWxezII0bOibBID/klQWUzEQtVkmuzrDmQFuq1b9QX7TZs0PhgdlhP6
ZJYf1Qs6lHdKODsy2uR8jBQOy0KIFe44cVUYx7VnafkcT0WZ8Xxb9+0y+Vl35xEFhxvC+78nzXSj
LNxmezK6PQwLP7VtrLzTv6ZSGyw/L+JGaviPZd5WfY/9bkFNVXDrJpN2LgWgHUCQkkJLZf18xeOO
w4A3hiRqgsSdujMTJDJ8s2y5no/Mnj9PWj/WSZLzWyzsxlHSlkKXFuQPub4KI6CGZlzt8/ReZo68
NaFsjyojDJerQ3w46lSgybLkpoozNEARkzshgstvKUq5LoF6bFntGpnuEUY19K+PdBQJ22DL9jcA
emu+YmSrgoUJgJo/vzPW8rA65/OvQdnYZiHQRM8VO7Hz/VD9dYJrObH/TZODGr2e6QcqXNo4awyp
hqh21QigoKuJvvLUStJZKVzjg6LN/h4xJUlhDWTsZ8/G1gf6pu+Sb/MhcFiFmL/VuYqo5JXkz1rl
EkyqbBCsicD0LlRmKXB1KsRCOV8rzFP1BbwzXd2ng4gY/FqiSHUSEo/4Wzg5ecNi19gTcQgEkI5P
Y/i0FYEXy2YYUkXtwTtHKjujQukABxqJIHBchSoSxswovcfkK5KVeiCHNJ/yKy5/Rd2mxkhWC+1w
9eZ6VdjlgiYlDbNo3e6kDTLGtGPZ5XC/09ifWbKrWcPLe4ABsbPM32RHNbsALvY0aNymow0MEkiY
Vwjgs6RjZEFE2JjMS7NT/YptlzbjeR5iLWu4UhuTZw7QhFsdnG/lamLa7Xq8FLXN70TZLDRhXElD
fYLUC/wHVcS3lFFvSwBzo8+XYQAJZcSWH661OAFg2Nuyth78RWi+HBbC60enF0ostyRl4c1YniZl
mxic0mV4KewI1ax1YGdma3h9B4yO+lcpNghVys5K8Q/x5/RiQRMMu59yzBdwgDkm5wY14mu57OFf
/RK7mIUqTu+kcGIxVZohxcmoNntT+PrkDZ8FLN6bsvF6mHML4eD47RglpyeLQ1VAiwTssDzNk5Dr
HFRIJH64mvxGADHy/Uj5lIXTc7SpVjFcd1NEuQKt/nmHrFedhagoqmH7RRmSrQ2Wzfy+IQexf9re
TIWtpmDCTl2sPC9Amr62so7nTAdojq6qgyrzlb4xq15Qxu0yVWm0nRlHL5sWu9gMdmEN6mIT7ZO5
bAoiX66IJu00psWRH34EyYRpGyHY0ChFXvdi0sWPHXPjBhb54ymrqsQywrjGsArb92i3e0yf6Aek
om8CppIhzKvEqUkVr1J1tQHwd21W8AQag/4NC5SMpcQCiS5F0PhTyIl1h+2fp6gp2vShZmDq1ODs
09Vpi+q94t5BeBPizn8BcAlPhljxKGDN8YPXGsBOPeC4oU6+7272ib3AGqqutCvVPXbGXvM1nul4
ZfqtWDKPqGJw/RnsPJ/lXUPF3Ehse3DQlSRM0FpmVuQAJ7aafyYqdV/TIKTVvG7TOlJjvNbXvs72
wZdTP2YdA+HvYd94DYjsgia2dX4KC3/eEJG52m8noYgLv8mJ1hiFb5X9nmV5vhfMd1SPU3fQOszS
ez8VEIWVcIO0yN7DAmo8uY3d1JBR/6iFO4ctthL9mA78eT/cgUMwa/7MJ0O67qJ95oy7dHc2KWvq
PW6PBPJY6SEl/wjCAyaVJZ56zJwyZQjUhbhBmDugI8kZETfN9Y6bcyA4KvKnGgbCstXNJe9CI5Th
kDmFNwUnzDKxZpo+0hw6uEGoqd3/vsyVi97CQqUfdVQZh4SQYz8E/YUHesETfhPesepUnVEzB1ad
LbGHtVG0dmxY0I9e1Hy9340DtwmvKlmPczFoCCe2Ul56ED4RI5hQreFyBieMwRWxedq81294Ucg5
EWgM6CfrzZFxisHauUPrto7nHlYsEUOJ05vi+fjOoPeDYN2C/xOf1D/cp/M3ZzgccCPxLlSulrLp
AXt6SSkV/TPPa6NjywyTyW8B76Ym5tezgxSxkQsJBfG6ABP2yGvTKbc2DUYEUSULfSCBhkYpTpae
GnrXuSILvSfExwRxXNSWL4oZw1zLInnIt7Z+6OKwN9F8HZ/ziLTkvKE5HYc71ZksEFSy1FSfYRVV
cdMwaMivd0aEcQoORtuY48XdT0MoGcMwfkK7XRKd5NTMbMqUV/zgVXKCwjCeUxt2D7yDU1ym7X5q
IiTzNV3WxxeTcNZObyj9nuiQQOF9q/Y/vMlKP2cnCjzKGRM4iFp6YuCLAnk+4lKChznltS66f17+
3AgGD27VqbfhpkdH631ldEBzH4HVC1hB2asNHrnjQnIpkNElJGaqcHLVy/WSUa9kzJBm1kFGQ7ZZ
80Wv7Tnn055rwvNvSVUBbq8TqupEDhboLC/8hV9/U7ueQhNm4+v0opGUkw2CyBBlj9Z8wn6Ad52j
hn97etWbfuKK+3YWmNZfVC737YJiR1p7I1ZKOS7+TfdYNnW82mIbKo5NYwnLrFfuAUjwM4LbWSqW
LZivg9z8ZmFEWB4BLPxxAZEWRqpddlnsA8shtltcPxxeA/shpqjsWb2qJO93gy2vw02ECkbbrtRH
nWMsl1Ztt8hgBLaNUg+UG/2W6uh/SRSFROgkQj/5pS45k/RuTof4om7slsSwLHtQl7F3r4qpzPE4
zZuq1+NPjTUXcQVqS18jCWkVPP38ZDmIy4fyGnyC4cy3Zu7xA6sXw0dy21lteIklfwSucEkVJR27
sW/neHB4A1aifG/9VqDfQ6Q9LnI3CpW20QCnLL3DZnNjknouQbbGZo9hqxhIyMvtaNeXGmG1xkXI
D3K1VSwypOpgOlaf2V3SHe5TPbYBoIagjE0wExsttTqGnBs6ZWpXX1GHv9wWVCla4nV87uVQYy3g
xNF0QSI+dp7G/RvakXtunHzsYShPkaElO+cN72/luEg5nvMF8hB5K0I/kzJrubmMYw5PRCJs6J/n
E15aClUPwwUIClOGtjmmmnfQ7tyQ5VkFlp61j1oOVXmF44WsXhwWKqgnjY+QpskmDzkHO1ELvUrQ
yBU2nkw1KYi5cF5CjiG27cwvnszSQjvqi8eIRPPT99Pye8g+6f8XFiGV/61TcGmR3MkSivYDP5nz
xK5BJEsUFFhgwT2uYO/bYRIDt5alC9uNrpDWY4jTcjaoXtSTrmAGt7Nyc8JVhKudviAy6hI1EWZj
kR+T/KahHR/8lUNZlBBVkodZVDnPiURN6w4QFphahX99TsQ8ufXheQEA6FFazrSG+/JFecukMC+d
Bxg5mA283u8h1TPaqLIjm1T2bZl3++nr1dfH8+zfagpWrQnP9KZ4Nw7ecmBwHxea4wORpAvVFo5k
MT0QNt+cf71tvKU/L2SCssr3dPr1rMnffpeoxe/JenF4BOvo0rlNv3hyFmt42L+ttriEeHMP0OfY
hMcTIM+vxVC3G5D6lfyBAgfqqkNvd0PNnwhhdqayyoAe7ZyBpt52jsIfwypOvvQSrKN/Kp5ZYweH
kxPKYY7j9GHBSxbeNIfzOQjC2olYjjr0Upn02oze/XS17Duesi8LQZKIVYboh9Dd7aKjWP1d9s+V
OzT4rs7QxFOJ3wNT2lduQEOwB0VIuuFRQ2ydxOeMXpc3n5ZiPM4SXzLe0qthm0LHXNBM8U8GRD95
xYJCJhi7PRZ1wdFq0yJL1NuZzHnd1RXmqAeHTTyV+qjSaw5OO/vZ4L3CCCIM56D4ZbaIJDwcbVbX
P6GQ9ac1BPUNSZt8EquM3VYOXcoz8j8SNTF8BqcY8n1teno93uPObtjCHdd9lYhhA+Tgu03s5aYZ
2BmBel45xFtKKWQXb+dxi9YUGjqgfs+9RCCRl+1uVS7l2XBN269tkk8zGAjybGIP4VOwwlOUsTFF
Ciq1qNNcbZgwcxNpC6U0Hr/VS/u7hiTm6+ycgI2a69kkVdcw5TJIO5+aVaA+hfYibZGfiui9DN8Q
6kI+Cf3VPkgznzsrHDcyFKl2LRxQ7DOkMY+jLchyXzffnoVEuefydu42E1dlMNMGJUXxjprRLujv
rolFnpwi771DwMFyAJgKKP3j6yblu5bU3mZvfM6hq8S3WBplBkxFSJOZvJocTFup0v5tmwnduvv7
kJY9wXzjngySSuBWEblZNzgCwIrAWkJf6FLqohGlACm+Y/ugj8yxYJ7HHn2UdTipyn2u1tNuEATS
0G79UmQuTYFv6UwkuplTRsOuBTOfieymUNsEBgzCH3clUgmlASm/6mba2hORP3psoJvedwtH27OU
yD0BTRHjVD5ICL5FPKEy7tzxHzDryARVREtmielPB8v7uJRJts6mxTblwKxAfaXah5v/Q09emiHv
F9g67u11ZmcL2UnajLtA0apJtdgiB0YEr/iCSn3VfdTBILwr4DrfmTXmmUMcM5GOiqDy5QDUj+dF
wJDc66A3fi/cxhmY1ZDpeOTJ3Iv/ihx1RxhgMKddKtgnId9iwqrHntLObGf81FohRIHmoiJqNr22
k4fb0LwNj2ntnq8TUxb8sl9A70j5cIVWiNu4rAWOgZx3sezkpUqgX6X16YpRZSCeqEFTD5yit1iq
i/a6FDp/ZubGY9N3m1VlbwNlp7DTy0VbW1JawRcvZ5RJNk2R1GcqLodIlJd5XtxM4dA8iZxiQnp2
73zZhu9ACQHJG1ai/r2t+F4Y/V5lfO2XLearH0HMZp9qwe16HtybJtudWFL9LMhaNgOL/kxwpWm+
5AYQfz6l6BtlW8kdWWUdJA0wG9/AfhjVryv0tt/ozsUsU71fgdPtKwOmsCe+uvYZkjY1YunaQOOU
M6JWfJ9+SLUOOC2mb0Y8DHk9f1/GrS05nZGXcyiwkybIGN0JGSmahmcif5JcY5kCLVSJEbhg+ump
hY+j3qBlAJia9kv8lPCkAwgNVxSbrafjfXmDLgHRqGae5fHAfvBnWZievowFNjWXtxq7zAq6x/YI
LZDRimIWOZJ3Ud2CE3Cq8cG7XFbAVZ7V9SEnulcKN5+H1X7qJ6fz42R7imhU4gfIiF/LYZRML6as
6Mh4mv7terLr2CKGfD2sMfS3PqRgl58r9qj6BSSL+U6m5Lfoi+vL1MZNlZiD58MFcT0BlcyblLCD
8YtY4KfrGg3PCpINzh5niivYO4ltaeBATUu/JinXvvswEkMWAvot3D30Z4+dPRIA9dnhahv4LZiA
ZeFW/1LKOK4upnB6+w9lzAH6tLyD4kZGjRAlZGuFmMX9eF6VVT+L7r7fkWHE3Utwuln0EzWjrmt5
cfte0OYFjAHyezpna0bDJsr2XjcD2cZv29gzDjAgXsW1CWU89MDZg1WSRz2UOLT3I6DqiGMdK+3w
9nWQbCQuQCUEuv71ZIwasr/lAOJg0HeMUfVH1Tms59yE7Qk358Z5gDhJC33W8WmUV4jDOb21l+rG
p6NyZqVNMo8lzarnOsKDHtdD1ptjFJqO+6djwQn3qPboCX33ylN2f7UeYwaOUGMuD6t7Z/WNP4H2
e1hp+shIpqTKM5QTfV0jCuCdaOTTMnMVtXJt7scXeowt66iotB94ZraxDZkd+XlwseSmUHCqBzip
zuvKbn1qKE4QeN+v052IuobVnyldkWhwYazq74svwBxwrLyVxGdEeaeH6LIzPJekUKJgulvbN8Ot
jch7AgHdH/Ok3diK6EVxEqSzKbRmEtF3H5FidkcZmZLBJNUigym9HV+NMkbzbVW+v7c6aJMvDX82
GCi9p7RNTYujxsWRLoUsqY6a16QpET0u1H98fqv52RguFTnO8D7ulBqds2qARqqEOZTWOFUm3Mie
+X5/CA9wgY/g9COSpKyrpw0zXrtxE2785Jhy/Vq1t4F5pHJM6Z9l7dKo8zpQsyVxfa+K6mbHO1zf
aWfqAoe599jvhMB7DX0PiZ1ZelZZJGNh94aPG44SzmusIrPgLBQAc6tuwBd29hnuYOtMdYQnlGsO
WguE8Vx//bKZNL+jBYtfBIpEXkKu4m3TuvunkYub61MmI68FjoFEYT7wArLuMPP0qHvjqRwDnW33
dBL4TMXtQsTGgGa0qnpYAe8RbHYC4H3MSxnLEZ9SZC84TUEK0nFobjhckpzP7Iy3hZyuPsuH5f5y
SLZgX/ERaRNa4kYk4kGfY8/7eXxTufiy4sYbLUFN9pivDtcbn1OhEMVX1nhns6Xf76XzvtzW/YE5
wHjtK+FHjgAHmBaqQHkvqYzG5qCU5Y91vDQROxh3IdWM/5UmROrf7P1wJa7tx75hdU970feoxVt2
19FDefU64i+IBda9AO11iYACpMQ1cKsvOlOFNHl7MirWhkh6Jr/J6IUisXKAXL+S4l+TJD2v1D+N
ob5YFsHo547LwCbN4/eP/RRyYku7Lw8fqyY8+Rg1XfTEeL39BjMY+FAQy4FgLzBHqnO62cada7Pr
oLInBSSVdhIQEvAazbOwGiZea0QVwtwv8wX6Ve3WqFeXq/Nz6PrKYlQCe2a50DPZIzOxqHELvg+R
fnlqcHS9sR/Mj/s1ZHNKaZHdbnOQXqE4cTwuraSNQFMHQUKlniyD9/5B+UVCJx2IGY12c13y0U9T
V29Jvz2iiXjwhcQgXzf+p26qFaEd+moyURh4ivgD1Yqhmjc+T+F1sP5V+GXHdnTvIH9tjSs2Z5ih
qL5THmctUSq6Sy2fpGrPO1Uu/qQK1bRWDpiV+kX3lQ47qR7s8unkn0X/b7Iry9dl+tUaEMOgtJwB
QeXOhHFJu+Ma/JivUsly9KCefo64JdWTujC8B6ukBiaixqjJacNXt72HWy4Wqs2W5dIgNRhqwBEM
FuEKnXYAG+J+OAENCdNm9Um+St5joixqY86HGgr3R8r2VKj8VbpiStyHbJY1Dl6+8j5i7T+FnXZp
eeX6pJJCXwbMITgZZMxLiHHmsPM1oukJ0uWt6Z8BZQpmf/GRkUCIHAYWODZBPpksGD6gUmS48QaO
nlpWRAJbkefbqicbjo/e6N+SzU7lKrx42JRkLFrWOinTrkN+pIEvMDauFiv7e1mRvhjT6ubE8F8a
8iZwnC9Ksw1PSprpcUalfOibudgBiS3AZh4j4HOaUAaJVWG4JaItjNr9PvEThp4Ygv88NU97LcHy
CaAOytOZmQ23L2mNHC+x9BHbyH8wPFUWds7WIUDDCgKwDM1i+3gGh51EVfbQ8i4p7VcIgFaLQ7oz
CLovU8GGq7T2rlEwtWye3JI84VZEyXn2znJBFHOodhI7BVJmexPuPIaaIKPadPO0/7OUp/+Qnw41
JsmWLCg+Ft3sv8ap55Y5yFA8rEBudcIH13q4qeySuJw3LPCV48fDXDeevorBhYmiR923Mb1KQnfe
fuC1AQpG5sWMKfb7XaH1BpNl7YstPKvoVxj8YMJx8TIgB4zHgfDi4petW3cyfx4OE/fgCu0JHAXl
zkhZchZCDFAB2iWUBOcu6ayBz8R2mJdmgHoYBQAIwblJ2hiOAAHuFTfbYwRfNIbsLo72nuaY5uCD
lUPfPuT7eLpvdl0cguW7NwlCPi8yaDw2t72LLL3nV5RjeiYxxFGl9oIc0MUp/8YlW2wYjGUifbMN
yfhVCkdxcEH3OBbOY2wZRXFiDOLTGXIMkxvfcOFDaBZaX6UHpkAODGLQBk5Om8Pwi82MRlgCQCNe
BcYY981xDUdE1DUkz4L/NRrphIAkNutU5thMVfuLhWjYW+NISe2pN9nRyRQ0EgYtE1M0OdOg57FL
2jsUA6ApfyRLkYt8ZBl+01JE8maw9BzvVmljKX/4yY8z8M0aCo6YUnrlfLQAqk7gF+jrBF+pt8LE
e8EmmAIXZP43dH6vhnc0/Qa5lXcKkJbwTHPbR+ynjxC6v6eRiTDsb1NsbEqsTEiTqWLcWueJG/Ki
IvR53V9+8IhuA0f4c0vm7vZ3Zlmom5iQaBBsEdefEV+ANu4Nlzr5p+jmsB6sFIFyP+StcJqHtY5y
/zueJ6JqY4BzH/qmEYTmcxauJmarcc3blhu/WeXlpcQQCybFroqux2PVySqsvxPm+A3AIHltm3Tg
H7oWXnh0ghEwT+VWGDTfCDCh/vIf43AeVWZWafuSVt6GzRdaA8tvw0dPk6LLQHNm2jHsEpgUw2zh
vwI5aOai1oqbugAvCqhY2XFkXFTvIGVPi9aFtfDwPJUIq76PP5b1pj3G3HsGZ28uwqXIS7DttCSB
TihWz9+WExINSy+E+DG94hLq8HL3HLygTmjXTLg9PkITDaEgewYt67K95AJix12DVFkcGuH8AsXR
IJIrIk0tRLjdVlRXLkDgP5lFvH53EM43IIreDH7FNM6iS+O5lIKBAG1F4s2hj++ve7rsd64CK/gh
D5ajawMgfy3D8Y+JBNdvqKCwMq1nyteLTja5z1mBIuaDFH8BlUTNVViKIM+exrpHJRCr0tJZ1w4I
GysL82kPRvyo3ZFWsd5WI0O687GUdmXHy8V9TEyud3UWUJpWBhIz9WpunRPokR37TmhtK5slzyB7
H24V4+q8aaFNJQZRJ/LZRsZWvpOVFgfmrLhqFWnQ7SRLD1TByMtjfivI7sc8psRVCibRUT7gzpBB
LwHcedKjEH6WG/zv6D86uDuEom5FklkDq0hIJOjAIZiaSLmCfQbRwePw7X/1vmHe39DjPYDtaXtp
A51TbFO9v1o3RCt2FjpbDGI5pnr5PRejBh4DviQQx4NUgbjU2SAYXB1mvGZTlfcZuilo/TSiDAyK
KHo+bsYg2c/uXh0NC/PI4HveivXz6pr4Otkywgmg/a5Fc6UqayYYQnH3A2hiOEwmBaR4vaoH9DpP
Aq61GSPCDWDMU26jv3rpWmArOmod/AU6zciW62kFH/ew0T/XS/Y4Auy980sONGKNSJsqyHcbboWF
LiizzFobBnR7z55vO1dcaDBUzz16YKYYUIB4cEUSdF4vSWKUu1kFrRCibUAM91BrsJ8DgMqr+3H3
/ZWauFkpIokdU5dJ1mF5nFvY6SK6IbgkP/SotuQamk3r3ijojTJ28zbJT1ZEe8ImOmh4jxukN4sL
nUEin0mp5exZckOS/Nif0iYF0dr5POP9k/CNTih25N3oHV5yaEEDRclMhoIOtHV5VPsig2kYLk1L
Il9Uy4WNKzqljpqy05ukT6ox+tk20f1Wr4u4fX/CnQ0xLgeC07rdJkao+5zll1RiXwnO+Enfhovh
mJcVFE0AATunzdxRAdq4wMX9AHTC0KYH+lCMjrNyWvoZtLHbps1+utDidfbMuQbFuBBsjvwR0Gem
E9hzmXMpZu+HJ7TrvZ2q5OqthlauczcA6WhIzqkwi/20o7Eqh+ubK7PVrqUPaz3nVxJ3N8WqD25U
Xyhyh51fFBK/27BfLkeWbuedwwI9uE6wBmgY0U2bL62zBO9au/FibPBU875ebqFpNA5xnQgMhBo/
OmEG38hlciQKWdYhp6mS4Wy6WXul+MsP1X+zpdCBP3zmAE0V8StgSLIlHy7g8D/Xhyn0oeLtDbJg
ds+9kmUurqgjVNmqo3w0Nml5h71B0/3ypCC5IoWSZJ9B9VULqI0O0QiUxUiy18BuasRbpJUPEVR6
3JeKNDlsh9Y+2OU5d6+gJBB0JNpV5J7HwqB6EgxezAVyOb/3ygtNUVz7W3PeH0fNYNT7h0vyDliz
+FCTbt5X+fNUu0Am/nGpr+WTBj1V4Sko49x73RXYMqO1xCvayWmRIYlaZ5PTMttG+nELmlWiEbJ+
LEY11JtwvkyR4DbYaDxBuS2njNmA8VlOE1YwYCaPeUcdaPmpCo3vflZQnqSVDscs7upGDXqODT6o
xD5i/oQ+EOwX9RBEgCPBTxeQlq5XoRsP93aGP+Ptf2Lg5b6Wmf9t4KpVBaJnA/3Hp9yM23oL66Zz
0odWvOW/jJXooyHnibWuv6Mnv/rh40iz1p0BwrFbzCPHcqfiW/QnP9gOUwdTS+Q4eZgsOjpXYstt
GV2efkoOIcxASmkDzWHM34inBeKqaA6Y1p3do3k/fKL8GtxxNYoW21n+FDYM/DkZ1EqJs8eD8304
G8IrTH6+bCydfIzvbnOzONJ85He19Q8H6sGIqNeMOWtJprD2z+vOtV3fHcddoC0CoGhfQBEZsDRW
lhW0okV95R+suH63RIaC4OQXjJuwTp8VYoJcS8pYWesGq2SQvmVMUgNRyoQXy5mJdOwrau/0Wwfx
9WTl5cS3QQFqhfDBbRjw5MiXefBVTFZuZ6r8WGG8dupZIdoofdobKPFiq8A3Q7GRy2+ivslHgkrq
NZiun9NJfsA59dqWBvaFQ9sy/pe1adHVFfPohLBYDZu/ucll0DBFRjpSBBWVzCYhF4jtsHPNh6jB
apH0o2kAagsEfb+lTGvjhHrYLlNWd70B3DsPPavvoic7jBqhqu8MulztzK6RrQjZgtolfPLvXkNl
Xezyc6rNFsB09bqujFrU1WDH1YXJzHMQXyS930a05Y7OjZ7OhDQLoBTDC3fSW2sQ4uvE1IJz2P6p
Zn5ImZ08P5sx33HHEc6G72pFrTqRSiHdUweyNN6kxuogoV11RjYhoXaKFNoTiB85zs9jm2vUnOuA
x1aK9l7akZzbzz2jb78Gmng6N/zU1Wt7RtqF0QpFzmkEshAjOnmo/k3dNKsbId7ZmVUY6175qBbX
Mm4KARI1kjXoqT6+llbHBLsOq7xvDdFugQdUyaCykJDqkrdVfsXxpbuCxV5Dp5pkz6X/ENuLgXhY
S9bHWB1HGWnws8OBcPlEaooVZbsaThLQKhx13WSkC2zT3Ds3N0AowMb56hE4exSpo3IrIQpUi6U8
dxnrmi0+C3SfiYLQKlFaY7M4gsoYFESgAISlWj5OdxyvFWTiQKkWhdVugB47Wx9yd/tRzi6BQP8S
K2teTKHVWUZSuyIL85reowLK+B0YGSoFyLNItKIgsCbPtllhTKc44H06o7iDsKRUI2OPVjTXdAJR
Xxuw4+cehn+ZrAKvjUL68KOZ34ke35EHr+EEz7yLf0HHw3zHUl2dTs7dPg70gsk+s9YsCxPd0S/x
7nWnFlX7e9GUtIw2f51j3TjESQmTa6V6qE70tScTERN0BroDRYvDyzgYoYALiGONxTkwG/uweFeP
rxooqyKclAhZrxnaNHxzk1TgzdIijnv2x7bV9X1spAe8l12BVPpjMaz1znvm139em00aMqG0bw0j
O/SoLrjUQmJVSqmL6KdF3xXmaD+8k+IXyYo2wtiEK1TR/xgGHpFbcO+jHg45JnABtlwObYCv8833
TQa803r4XdYdNmyuiFH8XIRWYjKA6cLft+JQqRd6SqbfdpZpxtJgANPUWsyY1Lu61lTOmVuJH7Ug
CjwjwPHPncp70gIV0K5FVOnfQaZSs2r9gsCHlHVQbJYBF/HpUGK+vthJCHtanuu8AoPX4s2QshWQ
SkAKpaRGPPeNA2t1wimHWHSe9PVmgz0Iw3r1EtQcOCnh/SagpIW3+B6JG9L7oDhNCfss7BO7yfkO
hZNCvDCq8qESa+5xbetgg3z0TY/pSxVRYBtbaPM1YZe9S0LxB4QE3Vhx84TQtwFm6bYjnUPdVxzH
3lbA2b3DVw0kPLVdWSIA+swCW8Zv1NtgcYkJfmQ8VtIKH0NIky+6lpzYLLQhr9JFEOCwYHaDis5A
2INrvJXE1BSyFFatC95Z2hwjA22suYOwRwlFVYlSyqHQiWdFS5xJ4k1xmHaUP4sKUmbQ91+GpSyz
YFNc3ucOgvipT9JlAExR0wPNr2YZ+WfoC11rZCjjVOIgiZUc8eJ3IgKSEuHTk2AyYvyjwVRSmljn
iR9YHo2cOR4IA0OEPAe0lEnmSfLdfcSVcyRM808vXDS2y6mwHXKZv27vU+awc+4piDZEbudWTsbU
a9DxK72XT9JlD2AH3OGDIuxBow1HFuqg06LKKWZK7xok8MkXEMKTasLf+u4KsQA5rlrwveLddzSL
wPsYM8AV/ZQ75MriUVD4Z+6zEdaoijpSDer4ZxGISjPzgrm/5lsrXS4cS7xJQnoYqV6PMSd0G2NP
GcVjdmQyoVUF5DdVcxVR4O2XkOR0aFoI77n7C7XTgu3RieEvrJnn1hDCXuecGG+JhV5QU/IFaJUd
PsaI1yqoLiHObFPrP2tIUAS9xh3NCK2m2Rr6fo2V6f5MKipjvcsuDCREtnNquBSaCiBrEkQAyZxb
PTWPHHLTkUaRG9too0MVTm47rGbd7oWMgXd4phbpvdTN+aARlWfnpq877HbbsBCC+I23OfWQ6IFm
5IkCX2zOfdOr8dB6R+Or/ZpP7+KVxcIQQ7vKwDA2blkNTNqMCgQUFqCRNruzYothyfTUjzsc8EZX
zCWRrUweFPjNrtPlZgGIMUccRRFS4GbgvFdm3/YvyGmRVL/Z614QIJy18jfXgc1pL+EiiHoWSwx1
LN/mrVpewcXklpcJRTmA/a26WEiFVNwD0aANRl9G6KTgmV19zu6uBWR9DxZssdul4AgAhwkdaXXr
saihOLHb/dsrFpvqf9G4iKGG23WWWixFLM6oMNR8GwushsAWK5nv3p9dNFX6oUhukKtW9GSO/lZg
lHSvhVZpHfd8+prYZ72j3sJK4/goCU1aFIY+M3+hGfzPLmOTW7iMAcXdYx2N0iMnzSAMs5Nz6frW
zncbebJeR4iAbJ8xEzgJLZTtcvF/lzI1AUenn9NExZm/K53JRNrqxm0TrC2fPHt/FDY1mwk5eIR5
d8UrNoeYDAxUFeWjTUaz1Vu6yW9RQvuvxooeBsniGH4rVO8jPh+/NuueuM3To9Go5mjOtMrrRjQd
HyI9MsFkEqAMNQNjtkfVcGwMAiALjnortfrC+owWbuvct2ZFjUZH9osbL4epogPS6tdCuKV5ABTQ
mGt+hmgghq3UhEkNH6Tbo4YkuKLZmO6nnfSAA6eKwZBeX9phSBclkXoUTvP07kiYBaBsD+xyQ6FX
xNfScOlvPlT/0ZAzFb3omNPzk1EqmvUuoBl3PIfGfvpn5P44my6l3H+iqT4NbmywXKOVnMma9Ovu
0dEb4M7vcFje4Ck4t8WirqLk0iZzcu7nuNv9RVA4WY3VOUYrW2UMy8p6UE93sZfwh2wObeA2fpMy
toAAg7Na3jmjtLcG2dg/Azo31tcdDnLLbjyRwAo9zyCq8p+lkFSSnb2Ajig4OC6nVeDuF6fNU+TY
BZX2pJt0g3ygoNzmtMRYDhRptaWdbz0OkIfdiW09rGJ25cV9norpFEaaiP/dGwV4TiLc5eubdEbn
cnI6YvDLb5UWIDQQaCTLXm/d4jX2dGvexKTEPqQnAKYFWh+BURLwE6fkmJaaDOJ6O5ANGKMgIGlS
PJnlAB++jqy1BtrZXbxreGNHlWtPDO7nyJy027AFvyGe8FFd9BQLoohY9oXcujdm+b3shE4KKnwm
L0XQ5VtXhpsOMKB7pWfaiKm6zCQRH9qoMKKyi468UaVipukNuHodCj6XmO3URB4P3eVfaUaCH9WX
283y4+FDkax/4n7zKeoxWoTd20J4saYj+8VE+V3ExSI56PNWcRVsJ9nUUjgRutMHxKpmBbSviDhv
rAqkhskHqxHhuWe4XahL2wEaSKZy4eVtLjXQBX010Pd9J3G93IVGG685scLHtGW5fX1XpadVW1me
PyIxLOB1bjXqr0vz+qd8lI2zAzrXML4iNSEw3NzzQWJw6O2VLGTFbThkDwVJqpg7ZzoYwjcezWXQ
PzRD7dL87r3GAR0Yd/ioRIL8nX7oUIeVO98DwhO6ihtsDSvkCkjulPrEq/VBuC3dJAMwNbEWmqF1
StEfeWUCMWxKOYCTXf0hFNj4cVCp/qBSazmC7lJVj6Cl8c9Vxh8jefJZp7ibarC9O/l1dHi665/a
a12JjYf+rr/bl8jXWMQbafBDberpcv4s2wWV0G/32NTF/rv7jzVUMw7ZJeQNyFZxQwYpOGBIDoQE
C9JFng0G25Mer6D46PKx8nvFv80ZV0RMLJm5OpmypwRMBll7r0/AZLgqJitZuMsCgaGUI6beHit2
gmycHD380JiOAx5AjU8cCFK4PI8PHw26QKybgp8BSh8G/4rIvOYGq0FCWiXc25RPo+IU+DonT9hO
Li83rwuFl1DEHOrWCt4N4ETE9dTaAFtJG2r3IHpGk8CroVX/Z14m4p5wtWEsdZUAlvU5it2KN7Xq
GbivledfnGJ41KDLxK6KM4JhybvrDMJRs3AVKTUbMkQ/aNzIGEAI56hTsORTu0cRQL21poFiFDfK
vG3dK8RJBfTiBxOoUNzR06DOYV97asKBaQNQ3sDxlnmzaxCuObbrpRrQEfl8+UXIseul6nWWCloP
R2LjDvemVn08SIIrQL4jGywFwkAWT1cCEdwGmgRz/8D28erU/x4v1IVKjDKf96Zk7dNZX89i38O9
ciU1UPSbCPJI9+JVIQEp3AFgjWoxPjcqkxB9ezdjh8l28dI9CMlIXOUya54T4ZmdW/PbawtGsNDI
QM3O4P9KoMaJGaJWEiuKUgB+lK01cnO2lnl6m7kf5nIyNc+kQGkKwqJDROWY3uvlxulSJeDoHYSE
XZ89N4yXJ+0EXuo+I0NAtCvEeg4aGRvl0bqWk4/l5+VvTSjehFBAkVos8A429XmT0UrsfZjyu9fV
zxd51l9Y18OehHinxVfo7zGwMiTS8xV41jIfl1iDch8akAqiF+bkqLdL/HUJdU2ZRkDJrExAvlFO
1gBfrkipJ6pNDxRn/84E/KaPYkXzklJRQZsTvN0zP1uIyvHsf+/n7ryMxdRY7T9gcixPkBbShG+3
324N9JB47SLk76+aG/qq3aVe5UQa4zNN1AnLJMXtwajqF6MsZ2dK7hq4u6A9oLpSQ4he9E9xIeOq
xzzYER3BK4k0xBq0oiwPz0o2YilfZcW6kq2SCRQDVfq+u9N7J1PcX5k3uAFVXQEJVV3dz5mq9CBl
pM3YhpDaYUM3Huh+f4dbLmocAVthwqcSM0DWhlLWrwM1KwDKk6ms1AystWds6/SD5NRpI/WFGfxk
RgWupkdfba1DxMZhVFVm5VPHYLtk5+C/2osxMu3jf7JS5u0eFOsN2Wc106vaQ2wcsC1DBhPOdDuW
brk2FccAr9Z6CFNdO5s3w9JDmjLDQjsEvd8QphPC7yifSGFbVWW6ijYFXvRj3xp82bxzYY3V67z+
APNz0MiJdGe/4pHqtKx1ZRyFzVz/fRBSACXODtC6+HLPd5AMmaICPC8bNLmMxGwd4CVytMatPqQM
EdRh1/J+98OTunWaEtnetcAuZ9fonPqyiqLVWWzhZ9DcfocL5Z9XjjAojiYqQEgnI7P8IDblC1tH
Ptj6z7NZLvLIUgrkwNX4T4D9twCDZ06/EMxc3v/LkEfa2nJ6QiYRp0IN1uwzMgmf8jri0XkRInqJ
pPtDW350gbJ7YBgo1q2oK//qNDX4DHhZMSi5DYUNrJ/1T1vYWng/4Cgkj0pSy7WqXiOBmbzJ4VRb
Uqv2tuDojLy/Ms2uoqzkj4yHe9xYQDNfy62dX3EkwffJoesloKESFVxRtjg4W8YFEuxrw3KFGkos
rlpFukPt521q9weRxpZ0AalmW8B39bXlb7wQspOdHgC/+TyEFez4RY0+/109vMz4d4ZIRa/ZmbPV
EmHmcTG58JgP2uzbS4pgjbHjzGP15ZvL+rdyzZGvcJ/PYw4hbiYlzTNVW5ERKF7TDGiVUPFXaZj4
kR392WXUnRE8fxyeDIT8ImW+vHGiNpahavbZZed96cWz13Z9UF2VoEKMn+lcs6It4z334K+vSOpF
eIVokoOLXydB2AbaMM5737ZgvBXT6b21/2+CtLqZIN9VNBQ/qT5sZ8JNmQLtOLqVtixONIQrbfnh
xr0I0NHfMgztEr86ECMLS8E62uy82bVECgSZcqeSpLqpSijpAAPjCVg+gB6ahqRDKmxcTECsiAJf
R63dyzGtJ62mlifOLhbJKWCUv6zaA4NWqAflWB6yqPMMEWtNVxhcKeRBFZx0XmBQJEue0t9KP3GK
1h3B9PJrdw6dmPLRjEd2zohph6OTungX4aUTFwlv4lUALOtLNMROwcoRxGs1rligfdpAUOYBywVv
mv8xUufexH0rIVVFfwA4a7v8/B6uP09b+XT2/1s3eenm/tBh/3AXkhPiZ8+oBuYeTlHVo/u/yFu7
mzvhYzHnCHIMI8TkVMsDdr0zK3WFke2OxgKp2X7X8rRDAcvld9IDPTOFDRunUsYb4xXIyl1ro/Y8
WiHRrhErmM3/rK1v63gxbL0itJQf/sQT/kr95yY/FRQRu9XrJWEVE1OndeeLYm2CzdpdsDM4BUjb
ru9S+h1i4JE+tbfjF8WBjSHWlRZzs022fhigpkQdiTMTNuRqpgxQPNpa9U6bAIs+940XiYpI9Eqs
4M+YO9wVk/AzuKh1b5XF2fJirjd4WJXPGxXtRDLhFd830BZaaL52nAiMrjKPtABYSCGtCNKgtSNJ
1w/zgkCKlx8N0l1bhyasUYyeYNwOaSDTU9CsjdL1QnyrxW010MeVwDStVlNCBEwra33LiSpKigAu
kA9fukZ0BgJ3OfRQRv9W3JbttAmdDW0Jjz2s+2MKLP0Aj9PwFV4nukICa5IYg2R2ZpQNnCaNIMQn
VcaHdCUitzd4O9J8DoTPGl1LfrA4qYVy4PHQo2iWSzMvaxt7Wm/rqUHI6BWX9Epsu8DsOiZNQ19k
PbHqGryjOfhlWPtCAXOf5H8xlLMY+tqzND5RsQItQUTbLFKD3gHMkscxNVqurPMYhSgsCQW0zTmN
UKPv6GdrWm8MwR7IBmS5p/kghG/dFK58fCzYb7aC2rsHDJsFKYrDmBdCB/DZn9hSpdy2MSIUUkZ9
vsebxFUtm+N8F1appnlBl3odhWXvjRiYO6AS9Ry4O2by7Sn0W7WmzLneDhG7ZXlVVOpPH8b6RIhI
QDb52KZFoi6pHIfE7AnGoaqIyJBNFgMre3kHOZcPygHAtb+X9K52/8OcWn16/n7zZ5+mmK97YQ4d
eZvuHV6vlMzpA7YEuu3fd7l27DI/UYO7tbb2sd5Gs/WkSgJSWGpw6khxblrSZt1H6LNibubcPqFS
uTVeFSuGRUjgezytednyZrg5PRRT+MvhXqVNG8FR+RuVJqkCOdCoFGlII0g4MUn10P9/IzvqpElC
AavThT/H01JOfW/jiTDkzuMKqhaO778C+WHzDCbJWj0gLHRinf7Rp/v7Ra7OLcHhUWVWrGToKlSU
PRa4k97hPwb6JvbUPD31jahw2M6MOCdyAabYSQsQ+SIhUMiHT/BHCRxwlbcZVFphpMsJiKa1VvHY
G+W4qwZKe19hmVSY3Xqo2a71YQcjSc41Iwyvv7fvIUPdLdZmagC2QVeog/r3qwiMenKzMQn/+aui
lYfQNUEKWL0esgBiuXxbCCOxFpFC+MASmYuZHG9HLDyv5DCaoSYSUBFNrXa4UUvVzRTHyX/5FQA5
sDOpz49aLf5R0LEsePMFc3t/L2ScU/ls8gy1/SurXgfkTq99oZID8ISJRmH7lpdqrVd7h/A8vwyY
xndynd6wEHRWI2TxOVoskn/eNdzSwx3foxNsFaPxojGCqFNiieiSdsizjolQk97AB4W6Bspw4ytN
eTEj/M31EYpMLSnLfctiey4xYPcuBzXpA4u4UhARmr7Sd+v5R0BHIPVxjtCDH/d4SQCr+zc90BZ2
ELCGFKFFGiYiqE+gj9xd9a2J2Ke1LgY8Jw+kgvWldRuOp5oTQtJO3g1U1nh7iF0uEEC9DoXwnYIC
vN11ecPUGIhPh/ahTf9aELAtQICku3OpEsHeoex/5KZymY4FeA+EoxIX/TIKQE35J7smI0nyLE9/
egmy4ghvtSdpnhIxX1Zm+IY8g+neANDYPAAE2V9CGV+/k4RNbsQcD62kgQdhmAJ5n1r+ZkUp1ISc
4KDrI4bw8Hd0PfomnjS/eW9Z49vYtyuyacPhs2k/3FcOIR2ChkyHrG/dG2A0eeB5BfzeD2T+gIhF
Te0/XPnm29byy1GSvragf2h6UOlzXW9OVtD9LKUrnGoilYQG9Q9Mtluw26kKA31LxhnDU470u22R
0FsXcFTSqtv9sJrSvxhHu+UkLBPiuBYxZGAhtzGiU7FIV1Uoljm6We4T7q0wdyEB9F0AkK+qJTX+
tqEioPGdJ8Un/7/k7E/J2GKoL7yQfuceP56Qb03MM8J52bVDNKjCVHs2wpPgY32lyjR7W9IQeL86
r3JqFwKJW/V6CXLj2AmcU41mvOH1QYq2mMrQs3zaS2DXO1Y21Qg2jSMImd2ZWKCPdgRb+MJvAquo
ZAgJpbkMQJvGqf0wyfA4XsPGCwrCy0MlLjfM/uV01ag7THfn7Sin4IUkoB5HJQB3fwrhyyg5Uf2u
RVeEpKZ2A6nyPbrPkCHn5kGwkjLQSMv3Q+bocQzcEo0PYh8CAUXLaVOEVRJiamkEzQn0QNK0arGU
5pCAgOwCabbXMfKVsyx3pDZFIenBvaDoFfd9kA1udsFl7XMKkeeYEvPznTERElOiGVHeqw7gep+U
0CG7J3aZS3jqD1p2UsXQpwZUImvfLeZ5VUo2Nx7F7KPtTSkbMqPl2tRr59Pv/hCdDt6FRh3I0LY8
5NsVFdwiiz5yaU39zyEgnPRrWIdye7P33uUo1BmBjvoGgTo+tSd2Tfihy3lHTSDXWOJrjSadQzso
DJrFG/3Ble8EgpHF21Mez+Zg7la8EI4w6+LXrnzBZZXrbdIf/dQZhc1z4A/7Hy2WueYVaXGVqnen
6orjkt8PHmtt3IcNTwagi6zY/t2kn6M1MoMarkdP3vYEQV1WBKJUyTsPjN0ZZzHdNmlcbT9Uv6yt
KqQ/a5z9nZoyIU2Sv07TUf1ujZo8cvDM+vsKW5fYZOXoH9M8vuZMPC93maSKBeQr8fh193W08VPd
nHaJiWp97ZzfLPsa/hbm7/3Szcm/AIVO7K3lu1g1O+kDDlWCh6TOmz2YLpW8sZYmiQNIitX9S9SA
vmalvT8Ytwp0NRDhLT0bg9v+HTdWYgzldvO0NiVqr8KkeU+nmbpTxHv2+n8NmyHc4fFeVpH8LfV2
bMNZ8buuGe9hb8ENkX5sPAmfviM4Naj2kYpuNS+bcH2UlwZvjHuUtqAn8vYulvvUcS4Mhqiw9alu
l5ZoazvRCOaHrshEt7v8greEuFEyfRKOfttw4kmexqc7DK9h0n+kkfpkMuHUzVUeWbW1oAz1U5s6
Ximv60A3oVSQdZ/2KMCXCCOejxKD2XcmG9nMZErBmH/t3Kok5iXqAA+nyaeHrAhwRlR74CUVMIiS
rY4xTr63efQSFf14VDqFghHTgx19iy9nd2deoIvt87tl8F3mD3x43dz0/DQg0Rnc/67pC252zC4U
qi/FQ+AmXB0Y3c5eyPMK4x5Aq1BJL57taIikaVtrN+gkxwA43RKxJhI0CGjjnGYM+WXlxIYFnxZh
G6nufZ11xQmFjEm7LhFON0nA+FInGW289F3NlUjTLWc4Fzm8Mjk6Rg+8azSAgzDYUI4ZybyzNrv5
f1f7Yxc9k6yC3YeJVxUCBhpSpe4YCS7ctvfYmKFvZlv/BL+IurpcztdiwsGSExkC2qF3R2o8uxQe
KZj1nBSGv4EMENu2B8w+JfpmSSnR9jOC1sjJvH2dOqWXHf/Pd6M+K+LQ45MbN0DAlGd11YXYL4Bp
VOYKFlOqSLx/LaQeJC2RtLa+9yT5H1R/B9dxFc9T+cTmUdvPFtDfEmdhd02mnaWrhbsIxW1cZ60A
X690mKLY02EPDgQZLrW/l0JWBIT0+DbN2cJXlUUI6WFcAwLAd5bRX/kVV8WJPR1mtXnk3cHXrFqB
ew3F014ais2aKj2lkuNpjCB3fSj68I8eui8bpZ+BhBeJx/fwX7i170g/nAxQX/eSx+UGbO7//xBE
SCZZMyQ8XCNjQBFyPqiLCMGu4pYrxpx4DPqiOtuCKTdiWxA3Yg5tXaMcJJlbl4ehfnv+zr/mF+30
7Sgt798rwTBuiFgdQr9ogjjewdE7UA8o0kgSYjd0qKkp9OGGPh6eZ0HWr6bEL6JcsAxaMHoZ0SyA
PzB7GYPWgaMLoSQsmyW+XdEN11SKaTyTdlpYg9IlAZ++g4EhbuaD1GS+VzZioUqfuM0Pp8nmaOYj
f9kU0kmFRKO8Q1e1YbSj3TxiVWDiEa4pG+hWK567El66zE9tX7xw+g3du6z4hBQLhIf9PiogDVfF
C1CZfXvu/59a987W7qA3Dqyre7h+r9xJm+HLuqcx4qISL+9EEZ5ZrBCOWknTa+ASxl/+BpsZX+D1
BW5Ze/r7EVSj3Y53qoSQixOcj/Wj8IVxYXr/YMNOIqY/oB7LC7nCC9V2Jq/i0C2XkpVDr6F4rcSK
r9cJrGh6ca6uMKk4qeosODERMil+bMmxV8iyIidwd6WfLUt9u2vyQNOzyoErgLVFRI2TiQItrWZa
K87ZDU2hkWjMJuEElzM8Uk5LXeAMIUNr43MOOAG+PXXDWRLw+YagAi+q9h8/osOPSzTSYvlEGc2Y
5jh/9C4dci5FY9GI4jB4BEcTnVe3HvrKxsh7Trn/oiC/9J/7EGB2JLndcqXTIz2UASGW0LtvCpMs
8NEBLf8hc8F+DpaA95acBUuUbmvTITuuiIixvxZ+Q+KyttcbK/hnRNev33ttAA1MyC4eqY8pECMO
HL78j013EuFmoEi8ysL31qZFNgy9SUTkVDlhrkMVeW4DQAzVvFcQcmh6ZIJ98lTNxKvo/AmXERns
0tjeKuSAz9QKfmEczNIlKhagpt9xj+kDAMuZn2uf3IxXJI7o0JVQlcUVIafdb7zeHto4V6WmL4R3
Z6fYZ2pTPJjlsEL+8zLQ38VUQs1CbyaQzIitLYVtEf7Cxl20KRxNss+0CQNpr5Swci9Zg90S/rJR
nor4D+vcIUn4Zy7u7gn/MpyaEelfoOHCflv7pQHUBpLaiD7G+6RIHfJvkCvt4iAJMxGSnH3vN5SJ
PCb0CwEOcSBd0krcbjjX96QuFxXonQjlwB6xofJJ2Po8QIGt1Ecmrqc54EbuvnppfMRz/rVzJyBH
HOWEi9tmmNhFEYRfwtGE8SxPphAxOm6ZIneiTtBEGJKBe5l8dtwq09xkJUzQpixCVdARLkYv+KrM
QkmVD/IXFnrYCYwV9htM9RlUGM3YIM4BsocaPbr12hGu78mKPCrmUraJaRejKthtnwPO0xzg2xfH
83i/9N0ZqDrmI4XwlaDHB0a/URKkVAi/2l2dQiIpqCT6MHcIplDaeJqT00Xymjjx3aZuT8Jm/z6N
ttRCD6vD9bG+uF6FR78L5b+iX4r/NFylT9DRzKdRkBwvYx0fbNQ4AhfWzhU/zFd3zg1jBUhuiRsN
fdZuJ/dMmIjwcXlu+yoXQ7+dAlb8EHGWJYudGO6f/pSUjPaXQBmDEZ2d8NuN/F1ph3In9Gil6cCn
Ap2cSbMnlxUxidT/yQ4dPWSfmX2DThTkGL3qxBcFkxX14N7GCHxxWc/SDPnpGvJEttWOZ8t6Usm3
RjKekynWnCbt078mSfeu+ERcbGxE1i3BVQPdS8FdsQyTIZJuFpcm2Su5he92DgYR/OL5b3Cmp31+
uDzfBLGQy28IXqlD14D5iTUycLu5/N9US+CFyZw+DPx/MI/e2mafigHgjCjlyzp4vsV+cZx7YHOk
1faxP7n36X1XNyzde/+0Pokqt5Jhx5+e97KZqpSujfWQKDtJOeW2SIu2G0pkql5xW9I87NeP7yqG
bAb6XOwRZ4OAKi0eh+lxntKM+rsaitcIX+XdPZSklgKZA7k4YaGm5b2VQyb+dEB9rn3t8LZxo3xJ
YIzoK3QEuT3xjCNA/DSxbWlfPQX5bYfVDM9vUoMdeYiMCW/RG+UA/k9ebHkFNe7cE0JAiUIHSmxc
ddkUprMaMMNCxEzbFBggyI47bXBgbN6Y8IJbacldGoF2nqfl3EL4+mX2Nu0y4hIPwe5pgsK1iIKK
xFjWpxRXVnNiQMjpGcLyZMywsC+LvCbQKkX3hP5CU8NSfjL+fY7Y28IwsSP6lmr+VD7HX05ouItU
DF3EcOlLuFkJMBv7RdqR+22eX5k3JzJWPzE6PWriCu51RJav5AihaXpLV/ToKthvOg/9Ha4JZFWK
bJ9Oz2HX8uAjX3B6dqkGMjrpy0XCquQQSY13X44YU4IQs2T56taCLQs4jL8W7TP4PUfrs61XxEda
MY0KGh+egLw1qvayHG53RD5iZRhao1ojYVDo3zvSPG/RYBPITCDkPFmNuZ4vz6Y1HFqlHeJvE968
uOuxtomCNg0EAQE2aNR9u4YlHOBRcI1ug3Rj/4cHJ0c+g4F3v55M6cHM55pVxC+iJ4xbbHZQKoFo
3p0ckzpiY+CtT3gSDxPY7P5poWyJWkhxWut2Ma9CQajVdaMRLC6XQQFHxMIcJCMMnOEWWkqLzz7T
5hgo+1ip4zrKJ1dOOcu/WbRYu0WmAKMxciH14Fc6Z77pEaQuPmrBegY8gH1KwM5c7X2xd93h36BA
kQC+uS/hzzDepoyTbOytcSrf3t8847jpAdzDI6yZAPLYeusRajt+foJYa4OpL20kpFxNsXhBgaAx
0631rhsfaHhlvgewbTB4YZwj8ozklGfNtdMagc7eLsVXA8/QZB5PyWspUCaiFvwQJNZ5r1w6DoLx
R/PYVbxRPdZj5vwyxekjMHDEREtPyfxCM1LuWzbRG3sS2XZeIxXIdOBb59U+W5ygittUTrvF4nso
voIOHLykPwCF/gvHUyjHwQDXOd0joKz1LIPcrcUGnkyBPvRseXbS36qIT6J3rUk5qhp63vITCmS0
PwJD2qFVn6cyTk7wn+wSoRY+0wkmJnnJ1TyJBRtJC6Oe9wMu0qkousobC8GBP30iTtostxVNwU3F
iBb/Vj7pSjCXEo4lparUoAM2ja9Hdyc7G/U2wWbqXx/RlPUU1SBty3+iLAgGnUJoZZ+LnqOJb1Be
DFgXg3f+oQ/Aq+aMhsCbE835gGSutIO0RT2fhVDtapxBU+gfqFQeAW2t/6S+jXdLS29wweG3YOWO
g/HeQ07uN5PrtCEEOZ2FYP8m/JvEvMzUARpA6iNhDNA9EmFlbLfpYjgj9uZJ/X/2S2xq8ckLkz5l
b/7unzAEPexZEUQR8J6tbZthCjOkVK3jaP4Fp+43C7VR6dB/JkZ3+3n84MrCk0jzYrV0IbEOo3S5
KCeUx+U+y30I1+c+zumF3KwbM7NwuFsHhE4+E1rrYA5T9EVPE8DH1WoHpiXsop++Jcp/iOf1Kq+H
wPjMOECHPHHeSoN3SIgYRXQ6EvBzSwC1GQzj5Cmfy1lHUXvtC8A7PMwa6mdH/07gEplKa4pWlk73
J+7ZUOHkIk+CF/YJcDNGKMue2GHtWE8XXeBT+hnd5zIzlqJNFdlDMYAHzA2B8WPQBEZfpPRBjyzf
KiHgcb9TVj1stGO3QA9ArEiL2jHjk8NVtIOGdqh/K/xsjSnW2dXWP4psiMBShD1DSMPKt2Cj+L5q
+FQOUQKz48Q0cppHDFzry9IQ8OsHsRjp+8BlTflGzn2+dbuNqxiKIDblONzTHRC4yvOJiuC5cGvg
avB7dvI3k7K0pm2zpOLSAZPmcnq0Wltb9tQH7q/C+4VTLulqdV0L2FrTh5OJp/bTApcterCiW6eh
m7qoCn7ykZzvhXt5gL5yTXSQLhQlg4cwEwU6OQd2kVGIz1StcXJ4tQzwJJ8i3FN79zjRkBGrME00
Cs3gnAPsrJ8RiU67XmyGa/mY14QM+MNz7rZRF1xtVTKX8/8UXA/P2zUn35X4Kuy8sa21Q1g8pfX5
bJffg+vvjbDqU9Pd8X8FpylmW3jqBqd80kalyENoZ2gmaREPM6b8e9wnZ11zW5QsR9wtjLLlGWV1
3A9whNzouMjFFpebOcIc3zqGd760x2ZYFLEfxOZCW0h+iKPV2M5BrLiQafz3VBApEEtdXNrLSKiK
gW236cRJqMObXPF7Cd4x2M/UrCulJHM0Ee0eYM2eMhXmO4Kx6R1hz7PPUurIc9679aS6+KAySJPM
E7OZqwnrkOuXdTZVGjGpwVX7pcoJY7OSads/xqE6tG7D4Ix6m6I2ALTzHSQO6FZgVijls0mBbe0y
iUhU4ZtmNLkBemtPOa7Ewm7TJLPxbon1EoT0GbjpsgN8BNsDJ5V4W2nVJPnjEzjYlCPTIKu7igHz
LTFoaf0WV/nCuuFmv49523GW4E/wHfOixiSqnixPaAn5kUVEoqDL+bFKpkdOWncapQFklKPH/s5l
dzvprrmgVuHQJWVJsX7jQfXmaDZEnZfBCe4sUr5Z4cE+wzARFn6QCVhAK9rOchJh5hpoT1vSB0dK
wCy83wl2NF4/OC9HECwgIUTKpqyqbXNVzNKYjX3ii8Yo4HiXYWLxUir3kU+jO5Biwe+GH0VdH5nd
QClewJ0D3EbQNytGo8ioJHn8VUQrnpyN5LrPsrNy46Jc4D6cWhenpV14DhlKzoUJhFXF3qmWybp+
3XXftqWYMF5534of/jd9OV11zVjAiAY9C9/F1WxKNVEyVeSz8C9Y1KCuZOE5FOX/BDga6Ndo2WGg
CJOB9UMXwb+Su/iLOuqOP8KfqM6qtCsMAXhkAUyhFrWFrMPpEc/Vs1/RBu0Rg7Qa8l6O7+DcQuXe
GcJQuboW6XrZz37bQSR2D1IFcXI7DDLZ2MYnIWzjQbQCZbtBvPQw4iflh7eIINGkR2/PxOGKIBOx
0Ybj+KuVYTCYoMmfcVkijA+1+6T+NiSykDevu4p98DhjpJjz74FokMLF31/Is8iae8yIE4p1jdGp
pPMFtWInL7S6cE6e3kq+pqkv2yNRR4N82/HKU8NhjWZn2UeF5JeSq5TdarB27DU22Vil8cQo2DlT
o3bimpllc0oUB/XDepXh7H7oCDcXlJZZ0qvFvnEjojeVYqvwHsyVPITx2JTEluQAiTmjNhOP+jqt
4Y3m7FltJPF4fDg34zxJP7Tr80aewAGVW2MABK9qoe5nF/LJXdJ/yopqS69DskBIqbfx9c1tEoKZ
89lWAQgSDMp+koyxbXl1DUSFa1b4fpv6jEFEbC90ZSQbYapb4UEh4ripCgejPe0NmmTS3MaIssgU
el8Uexyj14MzJbH7cAU8wDLjB4HT8efvwqci3XLq9hwbcblOSCh6NZ7Fh9dygKgcl8Y7HrPiCli3
g5bM8VeMZJFNcsDH+3epzW8QoaeEiTlmAcPK+/OLyZrsLtg/YGmo/zbIVA1lPBYXzVzHOVVMLN+M
RZWr+DJXAhuKTlYmqDU6uNZtUDrwhLb0mfrpnP6I3uJmBwvQ/vH9I0bHb5wWZ5JAtJn63N6UjETW
ABU0R9a2IbkrsaPagtT/WIOrsnW/NFezeRXvRdYYtHwyjdPdCOHbLsRARaB4cha1VZnAq+Ga+Yrz
1B3QBllqXy+elS8g5Jn2uC9bxZDiN6aMk5/P3uGBLEzX7kCQe8g1UmOAZjBoFFdMt+UwW/Nvztg+
Mut9HYv7dciWblMXwp8XrrTePkOZJOq/KIr2LbWD48rATpvQz9nlpRlRJDJpiQoP/dNYMl/zWYA2
cojYN65/KP2VYO1bccpnEHmEBVjiEXN2VB8HLsu/uATZvuzA9abRLwKZGHJJN0KfA2/To4NxHhIM
cFuYlnrose33fIB/ZX/TmEkqtHrm/qG14B2v8Op4h1PuVWoXBtAmU/0kcd735S+3UkCwddsMCwLl
iYZFokPN/p4pc6JgvXI7B8ZgjypTiFstdC/I9vavD2d8LucY37AGh8iIk25c8crVa6n8WD5TJ1WQ
i4tLAc1Toz5BulGpBPyebl5s0C1VNzhBhioawQEf/tZ9vnGRhWaA82BpyOsfEBRYSUYk2vCknCrC
nfBvLTRCkaK4/O8mcFXh0wmz2I2GGgTbL4GhKF/DFMyDpWH9PNjhJucSNOkX0EALER3bJDT4fdpe
wMnNXSMam7u8M6R9USdn6xZkTR2zy0nZwTM2DaOdjUfshUK8/qKUpk9RcAZamYUiD24CtR4VU9Ly
sV5wTXHPkKSWjztdIoey3OrND0UQ3sb9IG25Vfk8YwysN8OGbnC5OjWpNcnq7PhrKJ3qMlY4ieCz
xW7TxPpIPdYs0wDEilBRlzeaHhvUEcYhXOhn0jLj06wJ5Go436/l4NQnWUu4OozMqD4dJ5Ezbw/x
LMODIY+xW0fyXdciX1K9FKJhBxhJXnLffaGGceOEUeKxghM2dxUa34fiScEZGzZHRiZswqvm5/EE
btZnVm28ZAMdCA+bQ+K01KVTmI6C6hM8suHgOGjQbFHvFzpavTbWeLhp6mzHecOc277JTmTQlRc4
mJomODOi3CehF677mNwJwPcdzoXwo5pRs7qf2gxqAA6KaG1Er3WWCuHnUdzvQ70wXwiOeZdd6X2L
oxKiB6bPeg+kGtMZ/B6cGv7KtsC1YIoy2BHyQItFIFaLvaM7uquGL+dabeWLmONXEKmXZGyfyTAv
iZ+OouUpthsAz7PC5fx6UaMKN35kKxnpB7aosICjQUHSCgY2FnNZ8DUBLjZC2wo0MoMn1NP7E/A6
HvVhESD1oWHc/wX8iFY2A8gD8Bt1+2o8SF8UtvdURNwvsnWaNJf691YOmv4vcr9fyItTCVJownzx
PYXgQDKmNRKHfK4yY6F8lMQ46mB6o5H5iz5zFjl99TOuxJbDy1hpY9nthQI1ZrawsmvG2k9OxBDC
iIkLS8wA7F6CU1d212KQAxs3IkrwtH/HnfCgNKbQbbAIGCWib5NwwxoIykCOzzphxj8VjstDM6oT
nesWRQf9Cz48GyUG0nr8fDPNKFp7nRBm8mpqIhl0j70rpqKTuEALl/bi9MI1J/xevUhK+fxqjPq5
bfWUzQ3x05zPqaxvQqSWB6YZdSDWnSrkAmkCRsuNMagT4iTrAnASQFWPp3xONC12Ks7aoXQ9vm6S
KeVaKm7OPKFUh3fL6xJeUyIIBXqSzanbhiyKbkZsxbhq5isqtIt0S/nP+LQVQV14ZeElR9x6k9En
Ffbl+eFe1gY1659cTsBTKE/Kjqsi6rVuk6crMHReNEiMil0IvGHSM+mQp3jePQRESHDc5ghekrl5
f+5rntqcnyqQp1SXrtHu4DZXwbiWMe/mjovsV9axUZGx/oEXEJi7xiGH4ZLQbMVb1d/SFwaGo7oL
maqagUJte37IEu4vFakA/2eP1orNmxUdsVG7o++OGQcehjcv8lctrEhochBKNytbJQE7NujNLGQr
ovcA6/tDOU43OQFQl4ghOvoHB0KXxvTsKBI+5FtJoqFONzsV/qjvZxrdlueC0lsNcbv0KZklg/ik
rtr2NBVe8b5/323vWEihMYS4oEuL5beTxICkMrH3G0OzwrOCs9AjljEgyMmID71FHnxfq7Xd6yAx
clKtRWI+bCJBKSKbsDMAqIBPlLE+Ps81MH9i7ve6efx2aXfkbutK0BotZSVd00+/oD/WZqFvEi9r
Eq4KWIJaVVJcJnGVeK8s0DXwkiSoJQv2y2V0bO4u94rq6C1YdM8THUXK5bc9ABFAI0wuVlTkm2v1
feLMgfGh1vrtc1O3VOXpC8wUWhm9z2bFfHaH1pmP0u1D30p/HaDVqzMtFCMaC1oKZs0eRxSWDQm6
dviwDdSJ7qVBYpdujtJLVqba0Sm67p5SRYuqOKhOYy2HDH94ACpDDHFccUmchKb7MrVHT8Tkwn5O
IwtY0KohxhUcCKitKirPwm+Czlu949oJ6q3Oq5D6ox9IZrMEYuALI28jr/5eElQM5bWxC5AHJqZ/
OZeGnoDu8Yntz0R+0clHodTOr3N0i6XdgvVC/MzfREtlqxiVJyoMn4CkJbYCezT5EDGZcD2SH/Oh
aLlZ98SKuxzV4j+/HiNDqGloDryIOmTp4neir5RVOCSZHdceqeaZJs1n/ou9PhgWIWCRceHrkEU6
/RVZBdJe9hzIr9kIW3vfCXGX4NGhPvTX8X7k2tHwV+al9HsA78xgM2HvGO0kRVe33uumvuAX1Zcu
IrQ2+XGs6bhO3A5OPY6nQilnbYlxwamFD1RkHd8HOrxD7MFN1mKTbtFHgT6h4cdr4c3K7mnEi9Oj
ATPSn3dQb8gkIx8M9Zpb15EgjOXISa6sCGA1ZhWJdDWlXLdYNT3axNVQJl+oEbklXyewO09JEkPe
++874reUWoUUfu5XOQZjgDI3Q8066DKGPf3fgDQbLGpbkQ7QbNoUE6KparkfBs7aFWoMc96oZhcn
epWHp316oLY1TnanQrcsYgWWJg+fXTdhFG2LYGnGdvyQyie/PgIB7iRwMcPyV3Ukp/6gFO6WoHd3
mIz+fNxybUsXZFH2cu0mFblTtizhe8Jlf9KdhfuOAX4MqIQERESUtC6JE8zBJPJXbgjyKBEDUCsj
NjXDX67O0MIZcuQgXG+UqWr1hKiHKJoMoCTuy4hkROvDp9cS8AWEVzJjxlgc/PEhQ3/FVIzUtGH9
GZDq/CU1fxFG81FDRSd3uxXQsK3djHTyrI8n3UPXsXHhAbvISMmNxsVe9GjGP92hd/0hXJskiNFH
5zZnb/3UQTtc3oT5+PxV7EeXezamXsNOnZx2OQwhGSSJDj+z0+UJedQl6zKl+binGtyb5qmALw+j
N4WDFw+j3NNuS7nrOX/T5xiViN0RbqAdlZpy8rTkELj7o0eW8vaLfRpLC1ftn3aYq9xnvjFmXaAe
zbFjeOt4YwsQrPUAY+vpYIBcX4BDUs1pgleXZ3/MyrBhLu2pcepBX/0shaLcg2KMSHR/ENwViUHn
HEnjhSBjNN4vcVlSNyljUZHiHRIYJ6xqmGDghwJlWB2bs6HjLTNlTt1Aqk2nyaxn3p/bhYqDFXh7
C/hLeyJUzbTSE09x+1TK3STXJqdx9I2m6bSwDJr9ftI8w2aPiMtG3+RB29oMv/yGkHrhdF17YHI1
SFF22CryG+8Tl6JUeH54v2wRLUvDL4Uws31xUapHOIATc5rDpRF/RPudrrSasgTBCSOlMcYTtjNV
/j4pi4kjZD2Kyguzu8Wp06s6WJwn+StBnD/rKv7hoHbrQF8BJbIR4Aei3Fer6f270vWa6ML6Du77
dYgTB6Wp9HTQubzx5pfvOXYY+zX8EaSWJ6dytbSepIx3ikJWzWIOEFNXjZgWNR9hYJkugyI+VaTe
6u7pGZeEiUs4DuO3uGu/947aL45dflC0c5kL9sGir8is9tnoxjPDO1tzFvm9SicvVi7KrBogfZDb
RVAh0dTKoiVDh4HjH1CGuBkgme1XQVlbOTfzo2LaGQyF8DKdINRxdVBEw5eUxGR4WoIi/dSPrFcC
1/z/A2KaKOtJN53qnqg1IL3iJOc7mYDmgUZE/S/BMkK0zg7seRlfQv5mtg0nTDDbhn4/yTCR03r7
apm4Y/org9oLcy+kXxp6LPrs35tbhbEPpAjKEHGTxWLmKuLRLh+wxvo8ELENI9D7ebZQ3v0n0REE
HFEj0HpWVThWVdT9zvA8TKfEFd5qJoKyoAxXWiSi2faJ3NRHDX/5NCxNX2WjhcOMyjRyD6tNnzPV
kDblrUZTHZV01ZGldzK8S9bhn6EvQyvuhQlv4xHjyhEuctMVo4jFvnZT/aFbTNk3i64rzIxNOoIu
cPB5e/Gp9ee+pvdqBupC32SmOgHdkaKJY1W17PR+EHCznZmrQFtLGodcuFEREmkstU0+yvHggA0W
XLWDAkaz8tgsgvCIESRsyVx0kRX1yty2ZPkDUdgXuyT5hO7cDWq56JijeGtKn9jAS1gENo8AYdww
NDq4a8AagZlxxBkuldteANmrffOWHQGSmJFJL3qtLw5Wh8oRmmfln+ie5TiZNqg4N0gCiSGys1up
kJc6/E4qjxlevv85JDd1dBrRnpIFd+RQDlI+9cyAzqYhbazduc6Y4pq2USabg2UkRF1IDGgDR9sZ
0qgC7pcwa2JfXuLDrWS0CY2BJu4/FOtTK1A9ZhRj/gKDjtPdcFP15SNR0rv7F509Oi6QzLQ/iGKx
Q01FnWPlQ0dp3mGF9O4O8r6TpIz3u9MeCwWCV4x5LQOsxHc2IS1glJSaTfuoKbHMuqk6fC8rQqPI
AZdrMP5va4QfKbc1PxPCywUO/ZUZ8/B8AYDM5zG47hpCGO1LrXvuPWRSqc8abCQbLsEQCNyRNXdP
TR6dhhfqmdYvR0IqleIG73nA8zCUS5kcVIQ0WvuvGZOVA+erkELqqk56WQ8u8nEgGLLkoFl/1fJy
G9OKdAoStaJMxYrcL1YODQuPIJQN5+dDJs/1uCO0Z+kdzCyp3v6jDEIZJOfX2PXSDCbSjfOjD0YM
KFfUcxB7QsgLgPOaVNL/g4Oo2bQb1g1nuJMfdHnFv4nJ6ZOAFhi8EQrL9xxRNUUA+ZLNIrKp0HTU
rq40LcGpuwbK9qOPneRxFHkdJhUl1RD0XGi/1ZrmNgnsvpYL5Suiru7EpUhdTvwVegPMfdfU6oBc
fmyCPmxIRBKRmsE/xjHufSm1o+hBx8sjSVbYKjXlp+LG4y8KOrOVXtFZ5J0+6bWtQVeT+24P9/pF
rYwhNtHQu72/bBns6uU/337m2KSDh9bdyK0c4NTuSZXjyjeBkEbi5k34INBhRiNCk1QOS7iVMSU3
mEcN57WQwunj0p+WXK10NpavL7NV0VeoCw8uTHPfF6NDapaIESCheXhMk9zCFWrXaBhf+NoT7SW6
9meZzscBoGd7R8KPYc78XBNO8Q3+1HpuZlRE48OthmZp4y6EuNJ9Vd6F0AAEBr1clJXH8su1fLUE
10tJ2JdomvnMGcCM1262WEEo+gIgw9aT1ygcKi2RaPt3wFmQBCPuufQZi2won8MtKq10quta3A+w
NTKsjUsfmms2t4cBbaSJ6Q7nXjlzOWuI+V1RPPt1i/s9A8etIWPdabns82jiV/HGMGkbBobuaHe2
7CShAIfYpr1SH44oYIw3f1mRYd0nyBJ4ODjEZTBmYDHQDmo0FssQabcGytMWKVDpTqgO0nFzQLUZ
ZHjkCByvrwgI4je0nStNukMHHAJ3m/2hZW/TK+wSKYI6AzXMvDjfa+xm/m58jyfdKzx1SSu/b9y0
16d0P/hXKDNAhuo7VQA+kbtqZzT6JRbptNL+gGGjEQvfp+HK1cBJQcFoTlXeqN7Kpy9riiWNypvF
kP3ArPMgD0yrHub6VkbuREnhd+NZK0Fi5HhR1TALSvQyJm+47Z/oA/NQi1btQKwWVufzI6E6EBHG
fbL6VGxmYH940M2uJcrN331L8gplFTwWQfXy0ago/v0sR1SW6d6RjFsisRGbsW4DW8wYy7vurPFy
uNRI8TxxHs+GIf1q7aemMxSCt+/ut2sC9GOXhqD+eBPCGDZCXr5vW0Xoz0pp3k1uKb3pQzAr/qGc
KJo0Cy+mA31TSr/PVu74GyueO7fi0A7TtInVhyYhMS4gGHuLqbInxCNDkxI25ot/1EbgDwrNYKPi
yb+nx/F94ICU/SQnw8ZEpkGWckmQjDIIl1ITQeJSMl4tlnVE5XV5W9twLZiWThLruplUkmIxGFjj
OebulaOelAGs6LebJACrF3BaZvWIP7N+TV6c/ta0HAnM1XQIVIYx25sFL+rENX45wzoj9h+24MkG
3wum6VIDUGl/l4kFKS8lSQC18wh+yiRMj3RmSDPnTBgw/0Qvycva9tYWFTFARAjr875gkQSl0dO4
4XPpsglRaEhsaRIUrRK+21WwPKJD32YE96w1d5zqs4jvqz7DCgVktMZLYlbwA84mxoKtzxoK2yig
AkVWmFZSXWGr0MuoQY5T8RXZV8SeA+zUHNFc1djXQovx5lNtc5iK30c9xZb2JvuLbKYNhn2k5qpH
5yb2n1aM5srfYjpc8wZow7bT4V0zQUd6yYCSzRYEzYOtKTytKoxEI5eQ3qG4TUrtDQS3duknF6gy
KU+mzu+NQJVgrXi3NWb6Vp+VTx7y26s17XVl4jH7GQKzgwGKm38MMqjV9RvgoNIFyGAuXABFJQ84
WioYV/NSJa8q+sYjvLtr8XSozAH9PNipcJI9Lyi1rqTGzRYSzSQ+Zo6rxjOUT9aEgnDVIgUA1Z7j
KYFC94Dz6tfE6VEYrgtP8nCv5H1M0It23w0e/Bg8ZaURRp/uw3G2IZCIrT3hcTNrKuSrtPrHT+cV
bad1uPtcd6dacuUELe3oxCcoT5n47SHTNrYqgtSkGDdmDmS/TUHkHlYE9piSTJRoTtK3Hw0U8VfI
OsEvK+O+vA6tZxrQuwxKxXt0OeGwqDBntd+J3X2WSfsL9HnZ9cGjFKAZmvJgyplzVGA0fsKibF9a
QKnDCkr5RnF8TWVmtcLsLfxHuw35CMr7pxIMhllgWD1Yq6ehKdHBxqqVafZBIEu2SrrDCe4WFN1P
rIf7FkpqQoDth9TUc4rUT5FbPFPvknZtygKxHWeES4mztXMowLUfowr9jCzRTVL7yNbltnYcFv/U
1qU6s6YFvYJp8s8pM82i+UhShAJ9ERqLN8nXdqLbnw+PuOUGQXZxZHUWra+6pjOf+4Dm66leh6xK
DCAQZyShDyHNQuab6QKfnHaHCFhztmJ8yTN/XRwkeMTFXZtiun5kEwJ8F3lXOVjWxKNm/SXQF9Ge
3oubT6URlGg1q/nMy20ytBC4Hqn2j22Pa6tsFTbZUsxV0T8v4kBWnlisIKVYYJocQmQwmXRaqBis
AdwHYOU0wcxhKkO+lCezrZXncj/qLL+JmvDCLvjYjUzuaUZriCCgkWmWbfK26qMm9McQDs5qCXly
nPeNfFrNZWWnyVhGcTzH+e8/l44Hlsyb2Lkp41jzBIpLrNLuz0pKuKP3YjJdQ+a94P2sUab0mkR2
TXt/nGxZ3NrMSyOfYxD8HNKMAEqFaKCkcB/ixrUu9fGIlwbB0/TKUGvclMtIaS0lzKdqOxRkX46N
0PmiLpFDe+6JUqCzx2xalKF5rxWriyr0oV0MZ2sCrvuTxQFrV/WXv3bwIVzLQjccQ70kHM7eT0e5
vBTpvQ1bAmwX789ss7jsQ+bfDl1hdee03dP40fYFWkbEQb3YZEMgkFHJKf34hZQoGhsC9oYDlyzu
76YnXTLzV+3kqIUpMd4qlpscZ7cCp9FsWzVw3jpJU+IjCNtjpxtV6s23WfWXBHKpvhf3yxBRRP47
8dvG021yEuGewy8MWhfhyy9bNCq4F4jTnxN4qVWRsNg6Q62XUNpN8nOnMV0K5RunbsUuVMIYHk/R
sTBoZsqSacUq1eg2UVKnruPOOzcKEQDvMCQgpEDDIqKsfK3O6BZe0KJv6/2hP8NMfuRNsyBGWu5r
3PSVCPO1IxypDsDripVbx/POhZTPRUibdZ6YloblRetObjgCHbrSs20sk6+JKclIcbF3eVitd7rd
p6gSSphhL1ILb1ONa6UNCDr4jEiWNMHACvNYf5bDbfRpB0QJtA9V8Vlw7BuEQ7f5aCbqHggby9S0
+Hq7J26YCMA4anwL+y9PUVGgO0DFA6doWS5NDQ9DChgZcxYCL5PbP5dVwHcE44R5VWojG0T14bia
DE37IT9BbgraIM16+GP2Ve6ch7PlJv8Buxfg6bsFBFKazEcrOAhYEYsi79bjE+8vCHGRgWpuKGzp
3eHH1omc/byUhkrL7iBi949WlfKmSZkAJsD6aHwzB4VHslijgmU71dLcpK6PdcPuqTFkB89F1Y4n
pBp4Bcr+cq6Pu4s3jCpwmb5geVguaktUV/GTFFv03atuaec/aR4Hcy/UD+jdWO1mk1JRiph3bRf9
2t68sTD3M2SQu4GWvitqaSPm2bBL9jilIWy5MUxD5jjbQ3AipyFvbXN5PAJNrqGgTB8U/7AeucD5
jit3ZVx3462nuAvMHY9MRbyBakMstY7P6kI+v2Wr5cc18/qzAKax6KGugQu0Hl5kCiKoZDDCMTbA
Ua1anMWZU+2C/WyGpri4FthqOk1W8sViG0jDf9mQZGV9Y5UwhD1s0Lwd1udGSW1hDvAV1A7VFJZh
xhxto7jsc2W6vKQGsJMZ2BUuZ+E+ZIgx0kjdsNvhlpZPAjdSX3ahQ6vngfihAH2geTEjtBMb3lHa
tKGyureyOSQTmFcG8ov6ARKQ19EnKSXuuScJz1YTY+Xc6wPPlk4nlCh5gJOtBGoFy6a75apl2nM0
yUsPRK542NkfVaa7C/T7xuHA5ugL4GuuzNfM9CNUy4dSVLmp3dMmYm/bgyTLGCvocxZY81hHuKkc
MfW5MvHaxTiL6vZR3SD1Mut+rFrf0raGZVJhHeQFjsfHgUX3Q3eIPMbyYSEhehghi+aohS5aDHum
eMrQGvJjJcJQVKCNKZ3eCtbKyHri2QN0usJ3Y9sGQcpuqdEvVBlD7ksaq1WCyu73aQKhPjvAqtcj
pdq+Mx/Q0XfcPzzVqQ1lo4AOabPcuwfa9g9/pJ88QTM2wBcgw8uYM3nuGiJMpwDqYoPHrLEAlfyu
WBZ/ntvSlrrnXy+AInm3GIQIH5hmGJxC7b/JJgVO2Vb5cC6oxk/2un6ogEUCUpxMXHtkhywNCDi1
JuDLx0662JEzKmHWUH8nGhUMU1jtKd79NRs6sraiEoT2RZqXxDrDBXIxowGaRrxvrQhwchTxKZfn
7QAOh+N4Qaib2Yyfpy1CUEi/Np2hw4NUySRoZ6r7oDsvwJDWs+orCiHASJ+3MqHKV1d01bZIwod2
n1sCw6/wO7evKgEA65c2HrNPHvGulvr8yFreq3zdRUJNhp6+2faOfu+wONjWU247uJBOzJQQIPZj
74uk38Avp1uUC6nHz/fnEJFbczbrhTp07cuITMqduFVCbgBXgaF9Ghmz411nuux7ghtgg1tg4EZD
donMdWam6d/Q+PPFnZ126FgMWw3t2ubNZMsd9xH1h9MW0QK/lT/onXuf34fquLNvlsPBT9H8KH6k
g8mDRxJRhSN9s/EMFzmHBFSZ9Javc0cT7LXD8bNBX/53JedixOQC3AJPfsD/94YJr/AwbWvhSxW5
KOhleMVWcaTMmKCVpVPdaDLQZagS9+5LVI6HglzaihxdrLpltkPujlbAIcCAamtCf0sFrSODNemZ
QKKSLHMTuYnm5KlTIGXX6ETthH7jbHC7BDqVnO+sjnUvzO+JNLJ3dL9eowt4b7UkjN9IjIJAapQQ
L6qmkWB58Sv7BmCtCoG1Wh+r5+Ac2Ia9/X5E2zJ5sZkYSz1HtAlHQTPddi8hXSCsEDhAAK5OopJW
aSlTBB068SvtYvtYC+6Yekki2ORBxXS+78/gyVqVYtlBEIicuir5ahTe0qJklsmTP2YdOHn5HjFy
hpVrqdcq7qD+vcB/Panj6gqdTFGPlqTZXX3RDTkkJrqHBwPhbK7Jk9X6NdHkWPkV629VYkWTxtfh
Rh789vwN5AKRGzM0IW/2sKMPwTg2Re6FI03V0qaULoVZR1bZobMppWh8vbGzX0MSGmEkCQWpV6bI
2W48IoUhqTqxgrVXBDoaR2kPKpJ0b1QiVI1grB7SJU5A6VUCLf58u6WLga6LQOFDo4tlF0KI+9n+
w/964on6Q3uwoi4XXjNmfqDohX1Gk9vY4bX7z7LfZdIWhyhMa5tDtEuPrszFzI86ssy/UVCSDsQ9
WKMGVr0GQP/gIuYT4uiMM6VUeKpL51fqk8tt9v9k8nF/enaVAOFjvkB2qDVV325pc392BalQE/Nj
t5OfvA/cs1xpq/qLV8SOF/er9cK6YGp29Oza0PxM8Gn1xFB1f3eLXhB1k1XFlAY9m3o8b6W/Runn
k8T7nNAIh2FCqvtBbTEgrULQznasd/CRELapDgeNBCO9iZM+IdfrwfWK3WOVPr4pz8HSU8WJvSFq
zMma8DVbJ/+YjvycyHlfPZqiKFqNuRDcWDhMPT3LuHdZeM/BzdrjB15npo23ag8XkUisFlj7+yzU
MjghEB6d9CtUq8EWZ/C/7xBZYeMJA8xXpwBc2BMi7LNP2NowBOt8AJ/micoZcJGoOaIWEP2v5ERV
mzrwBKP5wkqrR/Zw/b9P3Q/h6g2fkh3wYqTVje/PvnFMkI01nCF/nooJ1/Y+OKlm2Bc7Lml93GY2
kVMVEP4cfZkF9LVicLKjbJdawhi628PHFGH/8AIqiaY8e3F9K35LTeXLB7DNiVvRfX8K9GoLZxVs
ze7oZU8w9fOWZwx0FCx99NAsn4nd+SdSxxKzxqUy8yAUOk+QZilT+aNL13cegATK6nNBD+wQKFR0
QWPtnRplG3JTCl48aE+d4hRDBa1FpdFd/oA46qfXqc5/Z7kw+ybAuAwxYfZQRB0PQk6TCguqbqep
644o+6u0hTdgAvi8r7yAM3vV+uu8NKVANee4b4MKAHoCi2FxaiFLEm9+au2PVNI6Taf7REdkbPy6
35GcaAfXAVd8ZnueT44/bbM+XI0+ha4tHlRk2kqWtfoz6JYPi1apbFGbGNRy1Mc7IGnArYpv8G7o
9xHlvjIaPKEqYKG74Hc6t88SJgl6BeFIZWAd+PHY9xZHHrWKsO2G6mpx/fj0ldmXmpJUcbmdg3lh
FC6/oHUtZ1t3zvD7tKMLVu4XbhntMVzZKyXMxyld9w9aHwWmWx2JPLeBda7Ewfzz4A2f+COwu8St
pAopS6bn+8kSsQhwnvxwKsDm/WDzAvC7fJrwgTE06jtAReBIIs1+jmxOp7UlcS+NTTJgnQcpdoAy
EW8T5GYKwiPGQk7KTQk2pLPVN63pHdpzkjtfC63fEa5zIcbMBSYt+xu9bkrxoLYAU1XZ3xBXAX77
Qj2x8EiH5ubD5LXoX4kJGiFEJAGksRvM7QBBUlLUPljjlOI2IcFU713L96Tsk66iagB+m1hE8KGK
MQU+OMLGXbuCmf8H1SsIWHdWW+R237CDEoguC1Pm54aFtjTGhvUEPzlaYgWGdV7iaCx4YJ7SdYYi
0wvEifizLyIlh0YdcMqiIutMQu8iZjz5aJGsa+xVSSKoMPZSNsUJoIgZacqibFCX2SoCIGctD5xB
PFGpS4L3Kuew/A/igLZBoWooxvNtRiDfcWAx+5/oscAs+5Ag4br/aC3R4Lt2CCU6DkSvDie38S8J
StNOCO1+gOOh3mlvTRbTydA/ID2dVxhayRWN+UQrChnzvUY31H4Fy0YOCYcLcmZB0EmzMkiCRinw
Xq2euf4Pki4BM6IO+lVGTIpHo2Q/Y1jEh62RJISvyQatYqVPAoiKCvqfRVr13FasNmq4o0cha/Qt
Gox6+1MyaQKxmtsmzYqrfwKwtDd+wfuSWDKYw9qVjqVVGig5c6osHcZh4b1lTKibdKVUUQbNotL8
CL1wdl4vr/iwpJj4E6lap88q5KXDuLOEuMwWuYaZT5qJjRez9oLWTG7quEavaOoy3v04GXweJy9K
wTK8dQsFEA0An+qLTUodJI/sFrMG6TJ0PCKMwc1T381eAguHxoErM3NfcuoDPuf1u+4EoC+Qcbek
3vRa7G5t0hPXozIa4VdNIbWWFj9z+P6DUGhXWkN/vYIycF71jrTmvMxCejXxOqSLaOSOY7ZohTl9
5lT0X7pGF3e4kZ+VTF15gkZDJOLflpiKR+ZUuCuxhSdlHG+djm5Jn92YTFPLtoLnyn3JzoEIsQob
Vi0K+1Wj+KvZwEhsZneVlLvNatvbpUpHjaRQKJqkl505JX3y6KQvU3I0SDeJEQbdA8uea/yhe9dV
zt3XpA6X2iKCqPxaNIPSQ38yBIs31CyxADDWtTI4wXuZ9CvW5kfMjj4wXr5V25lokiRupyBWteVb
eFqg8e1XRyrO3NUFL0ZJ1gQ6gLoMM3AVCyIyRotLyJLBsAPs8kU4lL3nxXHdmzhc+JLQDm2TFsFX
2BiBnbXACh1qwRyaUD6+6XOSBz3dv3UW8/gkhK7DBy/0+VFpBm1R3W2nFP2MEF+LIl+jcqLYgN22
es/AQbrcIchuQX+0h0aA+vh4dOPjBRKFvEBWOrnk9Qs630Y9eeV3l7xCZnBAzBSvH4jPIW+X8Xwu
YKg5+LOJ16g4oA252hamHnBHhAR7GaqYR4WX8bC1ZAWIkecaTr/bf/hAiYhWkpBjep0hEzRsImRs
6f3NGZe+XVM7IGaych2R1dUki6a9Z7FerMlGYrfHJSkob8E4ulCfT7THH5QbMqGI78XaO5dBoGKC
VSoqRdj+Nie0O2aOMA20IEBFdajApraq2TcVC94t9yFoVY/ivZi6/TSDy0N/T/sklEOCOFQu10Pe
o9M5ZIukI2v9zy8fRZUKn0LD1oUCZ/l152He42HlBeIBqcdgzJMlywdA379jh1m8udI+hQutDrza
ky8eVeyZiRej2pIYdrJKb1yM6p3D1KQUBDsPdm9glURQZZcIhrcPD/W+3OLuTw78hAscKGUMdxsv
uWNKJZNKc3y9+BvS2lX5UpezqOxStWXeqUFN/n7J24u3SWp9d8avOJhtUdp0M5GW8KJA+5Nj4SRP
pfcx/0r71XGBykUmti4hmhfs1tZgWP0WAZLIx/KLngBs6ftbxYBtnKl0nvxDrNkGa0ShewkxD2DR
CG9CkCVAcmrrhAShGdxdC/V6HMdYhxEHTRz5DEeZRn8HRCo77GGJM+kKbgttLEggp6EqzfaKbcWx
H4fTSjJSRKClHYYmR+5RIIQ1t9d6fO4seUeGEedND8Mjwbk9crj6xa5efZfRMjn3eVxhLwA+x4Ll
ecVyp8peDr635MRq+IP23EDcXzB7L/PwafTm6b+YFqL5jzP0p8LKrUGa1CEVFht6PHFFhQBS9LjK
XtImvAvyQgYw1dKRIwfAvfKDcnZMgGb3phqRVZlHRUie1c9r7eUqtoHVRF53Ko3W633dDywwLz/s
tN18CsDnaw/gENCwB8pDZ53yw4FYJVXBrhArT5rl7bnqmBwwIumjHmxYUa3k0zxSyoS+Ydcdpkr3
j/dtWl8wnbBQIUBGh29Zkv9INkUkwxqBSKA+aoKE+fn8/HkvvzET9RWhkQ8wCnAsqckT+x1d9Vxu
mqo/suxgXBIi2INgyFVr0MEVMiIt/yYkesPOZVSEbOildxWApCx8bQVAB6upD1mB23QT+Wvly8aa
Hr9wpUwSL2AdWQzMxEKSsCvJUm/uAb58Z89aVDKwT6LsTnY8urA/BFoX3W3ENlY0PcuOXcKmMvB2
ZTYgeSrW9FfjlNOPz+vyiTEheettK/HfH97QpfpXYXmCADd7TI4K+eXrgsWHcT4F5I4pShHP+qyI
6KszrGW4MN8NL+gQfJvjmD55/bYjToE6tNXiRAG8tkFB5dDwfdE/iqj9lHcOFUqIaDdKVuaKrK74
OW+zCxmGG2BsIqdZYaL8bJlUm65QZX6cRjGCGSoSj1Gz7z2mVRRXjMDww/Rygb09eLTdUsVztoSd
ODFMEGFrTXZC9J5tH0hj6p0RcGXvBTPK6wfctrHIbr1Q/iDuaHoptjcCruiGoxUsfGVM2+aHpkn6
FXldrA7PrO3BtVHUkAEuLj7VawBFrY23IckRBVGFsrmYbr88hWhXUQvR1IpkwotpR/bSDNo2usQ3
jJF5WDIs8V5hY7A+XAV5TWidE/Ljx164t9KehNfzLXhnW3vy6WSFKtFLdm/geNZ5sZWuRGCAZfY+
W98hNAG3CbzPqzhk3v0MKGKjb00MvBAEphfaH4tiPlXTjGIYYjWHchKrG+uZGJ1Ir1rudpkrbqf3
winQj2zFTn/qKPL78BUjUMZs4fc6OvPl0VAafOuXMPUDt1TK41QRG/NC8N61XMfKexu/bUZz0I7i
+yhO9zgvRf+WLevpV9X09SMBY5TSdtAJdAXdd9NrmfsS1UG9cp5allSaNGAMuZ0J+30H851dXQVf
bHTGOLnIldmAnLcayuQaDcMMD66WNxi00jM9KOmT0OPnTVRicAgQA11BJnpJ/vYxJqmgpy2Rhci0
7lvZ58Bu9zAZQDpVWqVg3S3Cc/xZin4hh+f1ONYqIqTdSRCrF1tjiCyDmLAWJyrwRAXtJDhGPiXt
hBzheRqbcDu+bNb3+CmGsNDKIKhzMqYdGXcP98D74Ql4ao3TeViVj65DVJYuVBlVwp22nArPo13N
zzrqDEiGU0ywqb14bNPcH5H+KggdvfYiZMXMkatzSKgJuqn4iwFU9AGfRSK032kirpucqnc5dG4Z
QjiLH0aAU3bghFhvw6wDh6/hYEtKfgYD6MgIfCGBXcXnHYAtLanTOxr8ExYwiqZxqUO5iaVLLaBG
X48qk4VJpfxNu9bungVhiV5mz2UAXI0gZDMOqH7WnBn5FwGijtLqEviMhi/IJLJL5rogDrfzGMAS
eo+tbDkViB/m4x1EfEfQoDdu25JATuv/Qi/Lcp0XksWTRldWI0YoNQ9F3IeXNfntHr8DzMezmJYx
alBr4DvFqsV3sO+cfhoHrEBNuIm5vjcECfBvMhHepFh2fEk4rl9vXo+fkGYcMBgd41/WMtdMgSY0
z/9SWco5vM/PpqEY5+EHQwEzWYZxOMi5LzH+arl/6zly6ofbj/ayEkkmi0OQ8SL7gtwJcWWUtC57
q8ohCvc4IkA7II4PSe/JX3wSaUJccwVSjUYiBIdXrz1aiikF3MGeQ0Vi4cbh2kC+o0kv50NlycOx
3upVyYIqNeywJ7N0XhzGFr2iaPwjlMgyCRIrn+35l/ydGK9rs8gCxC1XFDlluZqdNFayKRjH9MKq
/wiDKlIO0clsGpWg07KlygzksnIXgIdIyKcTqkuHxfAYrslMdX2u08lTj/G4fA0+bvFvN8vWX9Gl
rYZxceJnTsMUiuE21WsJ7weTrxtTzxSxboF/wEyIq91n/mepqJv6mz/WKogXeaa2qRh4tysVcS/0
fsOrH1Gj+vB9ST/L4hrbqrNo9M8pr/RkwhA7tBNkboJPf8/Pey2CrUUpIQkhLNP/UC2XPlGYCGdU
//eKjiww7Bpe02qwfeNHDZYdSq7LZcF0c1SFXU4vG9myD3EN8UjqoD/i60C/gPKxiLgKKJXLi/f5
8ADsE/AHkTvPGKAyW7Yc6LWK8d1jvYowCAqMhOx2p3HTMi/E9x8Pk2XnexfQCf5BIBea74E8u0K6
ltjxy4fMg2YgucpMIVTx9clcFQktlzpSYz+UG0sUcKbGDa3STIcqCMFK8HlzKk6IhoTfH4KBCBkd
VqK2xGbEpJqC/qUKrD305v1Wp9Sst7ndAwdWyB4TLErdqqKoMqdQ7yhZuTPSU3XPXtfvDUQ7yWhi
iSOQ9Na8JcqVEMsgVS64VUWz0BtpkiP8OnowPpP9oousMi2pajpEL4W4t23RlT7xxiJQ+g2V9nJ5
vd116OSVcHleE1eTkFnut3FjAKkqYUprTc4Ja8vYLbJeZfvbp+2ebGR8RpCCRh9zSk6XKWDDZYdg
n7c6uyp6/W8ls+Cfx/TTUOSYOhrnIqVze3JbwlxQW4WdOIsrozrbMmEJCKQ01kp/GSiC1mSzBdsg
MDvVLs8ghrW+U+yCwuu8ePxkpimXnqbmjaZ5sslIiV9Zo1Qxtx5/+hWlsP4lrUCZY8jbf1s7mnbl
ZAYUG1I2faCiW7yuMFWknElD3cT0Na4mx76Xcor0xGQrfo1ctWiibbjYTCvEi3mTBIE5KYZTK03q
mCBc/hf0xTJ1bqAj6TJCeoynb3YPx3eQSZiXw43UF55UnK6vj3xacwtvRUrbphHQOs6TIF5ntgF1
E0j6b3uhkr2AJEp/AEuxsiiS0XxPYt2+5IpTrTJiz5ij1JULVOB7V0d2X3NP6iDWWULIQvEPM7Z2
Un4oXGQcsHCXW5kFWzgo6MI2HQZB0c/1wP4IKqNBrfcNu4PCIvLkfT4At5ULRuSJfX3nrM6t+TRv
HZfGPlOh1HxMrzbBr4aQ6TnBR+eCi94g6iOD0Kroej88HtpBnYeNGMR2qc0H8Vgjl8yHZLitk7GR
ACQzO6r+T20RzK9/t6TtH5Akuq3oOGB5yKCzUtN9pn0atYdShVTqgFTFZklbR7U7+hUaNNJySbGI
4GlX185y9HbHEGt32yspzuZL28txrUCQyfFcAK4w7oPM8j3+Op8xolvgSBuoIw4L7wxgALDsDiIr
UIyFRgjxKoiceYKEsuxyrtnej7P+TCEuDZ891Q/ELT7LhtTHi08haosKz+Ff8XfcEILJD+PooplC
NO8mY7mZxcBtyc8xop5nvV2vbwxgwEepJQWq7+PqO+d9SL+TkYCCa8EWD4crU05NRNY/52o65nTZ
5/jQz0rQwCa7y8q/Cr9szArL1+Xa0nIDtFFLx5lZiOUdOYF8ITmqHWf9Zjpi7DOTl+wHeAogqsbt
PpaxwrAzDQc32gJwgls/EZjPaFP2HCrFcxvtzpcY6XEJzkxCk+ltpmaX/Bk3ch1zvEMu+UOVYKO5
jTtmaddh0q4zIOxpCkD5QMZcWDFJFpi0Vhp8b9NFkx7r2zF9e6i9cwNVGlh1xW8/JsParced1j06
P+0OfXF2ay5ri8j4JoPQtzPvV6y7vL64VsucBVMy1YDtVT5KY1Xrxgq9NV6qCcJ/YtO0rPOZRKat
dV0mAGZAN19qtQzLYFUsA7gj99pL3mOdzzLsvtqfZld8bzSmpycyV/CXPqYp57t5QnE8V6pg869p
aK136v3dzovY0YA/OEsQcum6vWQpFbUrkH5oD5/3ffPmSAiqNYpdbzWPHFaKhjjVpk4fE1Ofh38P
NyRHlvFlKugTe3CT9KAFsvvk8bQ43GX2h1qDuIvIsjWXMbQ2KtAJffCjGfsOzo8I+pAnWws1Zhst
HS8QKE5YMXAAEQdSkkAwsLu5qEZ8g7pj6Lm19TlqBQYutyuEw7je9Ldo9ygMXZVcJJYtFdsc2HRX
TVBDd/FXSuXCtphygXg8YtMc5P+bfKpWvWNN5FdeBs3Iwm97N7izPVZV4CmDCFMgqH79ifVXmp6Y
eV5gjMeje5wpJNU015uVAVymzf0gRGlsEbIhIlR6TJpMTWYno1ULFuDAim6zkeyYYJnrBxYIJR0B
unMZDJ8hk6PxHbUABKG6sYcO/SKhwUlhBiWLZmKxNg5K++EzZtKxmOnhntLMcXWiu4STOc0WGLcS
Prk+2Cgdbh7r05gcN2GvGEfFwytiwMvAE0Zs+7Ayze2ozSi1C7C/zVS7hnEiYJgn1OqSaFapB9wa
KFzRKdANDdwmz1+ryNDYk2NxfdweYX9891+hJBc5f52i/c/gGpyyJmSiOfPDIoWsKHhoMm/wiLJ4
Wc2YSjKXKsWKyMtPLnZ6+p1AmpJYLipN5xs5FQRKipEQkZmRa16KbYhuPm/LiJhSPipjhvMtHFf8
fGdOSIljrcFuC870fNw94AS5QD04/80RulcOD2w0qz+F2Ds8QkEn/ZoRK2t8yA6ONS981VIb2pJQ
ZRNDZyrvvSLUI5kj7e0vwo0GgPVnjADthLYFdTWMVespCJOdePfMn85rqfDOF0w6pfS8oyQnj5wO
AsKvgc6nzNQC3JrgCpdW7EKLPL9muVKC5kf07dILt4VVh80+7/RGqRdrL/sI9DFqiz7eanylYZ7d
5AZHRQR6VgmdvdyD8KOsMvgIUGYX0MtAcBEgYpA2NLmYZWfSS3TIYtq1Gox24YctpJJdNVfzlOoi
14KDcXFkbtOe5NihvWfJnpnX+nQlLGQG+oXjoIxLJk8zuDt+kSNW5YkiL7iGvSghdnFt3lZbb6LC
QzuRlz2UB8ekxi5YP21DzQSZr4VUJwBziXqyTn5y+1VHUf1a8AvHAgwM9Ai3cvafoB6HU86hulPm
YiXC6mRpD+BRAU5UZoZfxzVxE+dUTt8Jx/s5kZo2PILFzXeiYSnGsJQqpEdy+w3vHZsCmwJmK88x
4h5+tPFljgX2+A0K6zr6CqXnmazEfUydeoH3t8cNqQG1LvorPlpaWwgaYZrddpaZ60Xmvc7UWClb
NLT4A9vWKDDx/yABZceojnwGFgVPBgjb8pZxXLZ+MVQ9xq4/E3r/5ePLb3zqH8aehALJclkZ203L
E5wZ5xQeM4A1Q9XtzwIgvu+icCp/SqfLaShaDvbwuT94qX5kdDGi/RFiyBJItzw6GEM4mQSpAbga
dQ/YterWNSyb0n0Q03K6jh4lOLCYRpIrq0jsPciqEPVYJTqgVD6sdapLcj6FkBqZUBDqlOP5k+XE
OPI4Vfo1clAOdpBkq+kbEdmRylL4TTn09/lM2147CJ/Pbo5NRf7SapZll6nBs/pgnEX93JzJIRRx
sSNWsDymqlac0ilFVJPOtRZ9FWKPKu5enT+ydYvA0axxV8qkuf5qZvBlw0ec7u0yFqopnuHPV97k
cI14BYbphLA+21vsP56fsYQebguN14qm7QOG0zBu2szQZXVW+3tT2C6j1DIUFsvGSPzah70AoVSc
OlARU/PCppOreO7HTaaNItyOSKc5N5jFj7/uTCOypH7UyG4yWz/z2T7pedoRBRKD44fwRCeErL94
bv4XElKtjZy15Hang+BO4l2zr7C5uyQSiTYwEmrxhHrbGhVOaez5S/CX6CODI5gRJ1HiZXDX/x/m
k2ixQhVI20kVHJoXKO8F3TfpgN6SF+Z8XoiFHJsGzxD8s4om5Tfk9GKGQOGlMMCkK5VazgRUupuT
WnH+Y4vMcfpAorR67Yw/GhtbxLCMtzB8oKX2xGUym+Gtl/LDZlCef5ATOgOchAgl1ivepJame/2d
nZt5fv5BUEEt9fQ1q7z2xKxL5OKmFcGCApIwwvJ77LRcOyBJq1gwQuPFqnOuKsb/3R7kBiAvwJqu
5xojiVjY5BWF7Dm/I9TGw0WvgL8aTVmtSPpgdORU9tQoIVKVwC9xWMfC+PHuGnNOp2YKd6nzdrEN
C/3rKDA0RX/VUmc1BTh34eDpXXeDIb8kqwMzXvrEbirfjqp/SzVxDnEtC86E5KeKI4i+zvx3ZELN
R8+gJikm6bdTmsFlZwOjYxzwBSdtq17byS6QB5nmo2K6wzVsz5e3R/68XQt5MFMXhX1nZtX3gNEd
Xe2ku27TYilJUr6ZenPlOFgPbdNfqcRRmx3URr06mU2nb348XfHFy4U/fRsMztl5OTg68hKZ3CCN
T39fBWPokPbLmXTN4u4PmLCEpB01fUZfmyq9SHhrf+IMy1jX08gegXWunEs6mDPv4QK8u2AvVlkE
SkC8ajhG2imAXFP7CQO1O2gk2lx5/yDjZCe5iEH75ZkNcRLneuonDbxtx4PPbXGaH+xTA0fbj+n1
WMcdE/5eC1GB8hjfr84vbmIYdNIVVOqrduvLTWmisAcWKDgHXNNZeptClHzVnkCaC+CusVRlogka
IOKgiRfIU3ECd7lQiPSbGM3J8MJlUF4n6v8sr9dSTTHnjgYeT1B9aAs7SjgZ3jdoTTOF4rKnTgjK
OcSW+qR4TyXdpjbcpCwsYCzaRRMjTh5BsUrWs0Dz78UDOUWE1Mg2MHkUkP/N7PtHAG7mvCuoliGY
pkDOciem6LmEbCSMUEPx7eaV18CHCU2mmZNddGXm18NizisXcnPy64fPCqXCg6YOKhrab2S0Bc4O
t0+1UP7M/dTZis/yllntbVBwLPezPJeZHn7jhQsysHc0l5ccrFUi1FWEKzF9h0q1b4NFwwDVH23m
X3QtymFf0um0PzkIr6M/qtOlX7xtK3pSVD5UE7MJaj9SG7IATwfJS1zNEU58hidqgk0gCCBnXWFo
PgbOEpT5LzihfrVco7MVtloh/+QzTHf/MLGY3cvVIQpSez9FNHMXAKN5ZPnfkGJj686i0RDuXwBI
D3AfDZRWhpOCWeDawxEFfZ911pXv0RzywRUWuu1Y+yJnbWVeZSy1qR/XQLFhmKG82dGHb7eMHGKb
f6OCsnGWIDLyKYq5RJNU6KJkUxFNBBiAHPi/vvHs1S/9ghBOwpOKWgl8RiiYfjhATypP5PKzdvcX
3KadXVfl0uPekPJF0KfzoNJxAXcKylCUY3QuhTCq0EmmOO6gE5VMXkYR0cn8646n08faf3xBikuR
3ncKMP0kN+XT4+SMXUXGOQVNIoTZ75ukTGYOpVet5IGwa6bO7WK6DApTr1VMjZacqMn/3lc2fKYM
VSsqascdFdadbRP5Mh8XDLx07pGY9RcEZV1YerhljoFCMIUScEyEXRaku1reFDCr2L90vhN+6rLL
ADObSeRFnyw6HdvGGELvpXQmuDa4rGERbq2j675xc760RyrgkFhbNmjT4Lgr4PXwU3xq3asPTCEy
r5dMVMMYf/KHp/Z5+Q0/Ez7QeIbAS/wFuatb1mOkye/PltHZUuRuIKTynDll0QQZHxwaF3BmRWWb
8ZGiiJ5jLHBfWqiYWTdqjF90dS+gUl9Ogm56UKtuT/aCmN2Wl1MalvQCaBeKLrji8ZwCpNrAsHZg
9w1bEcEsm+bHTUQlwlWHmEKI7rPcIEQ8umJwtQwSMK6uTJziXFWNk3Zuyt7NvfXNKLaf0UzgTYGU
35fQdS+3fUDoYKevrk9XWwNqAHguBWIkX7py3Pm00Ad8N/ruma+exXnC/wokiECQeNRj6ZaFkyaR
yHIRRV9y/0LsgMFluLj6kOp7ybujOCaeylkwBEzT/HVULP14dXqGvQkuSM8aZ4pGmIXjco/ksd9z
cQqty1ucJ1HAfR914a8PlZFgng7NQjZeAV0kozuQR3pKScgfJk3gmJ3Eb6lznmwHdEat7bzFJYzg
Sg7BnNARpidqyGGpBwy7MDNc55/LQOV4JQmsUWIpPaxx/NGld82NUxlTP4lwGoNbgfB3QN2/nifX
IUlwZWH7tQEFqS0RZ7ZbyPGKLP+u6VkFnZP4VsMNaan7iVacV9QKKMdxq13B04rvDIZvpNWOLIOQ
8dQP0xRj9XqgJ4uUONTT5IrM4I2vKXB3/kMzxPZ70d3GkvuV6c8hBz9s50+EPV2HSYDJVyIabST0
acr5Q4lIF/WZVjaoIFE30/YgD9R1ZcrYQR0tcHgEffgoEg33ivFH9P5XMoecBr6ygSSgRQSQMkgk
ZNEoEgf5kgWTiOinH/Itzgy0EO/7JpxDjKAC+LnkJr6x34TEdsl+j90c2OZdwM77Z7FwfZUPkJrD
uSLa51GZaB9MMz7inODHZ7aDNTvZqphvn+eDoZkdDJR6fwED+XPX659uS3OUb3Rc2SsxJkS/TQV9
bNGLHccqxTysDcJnfM86DtYA5VFFfkXjPQdbA6gqSrnb/+vDjj6tSUsoP734lMtBUL8eIqU0kxiq
EHagH/AAtmykQesar3JBA/X1+ClKga8Mir24M2N8rWnVsST55FyDPmV+xbunwhC4CzQhinkUhaGX
fit8kEum2ggtYdeqt6As9wzbaontGpKemf58E61kfStZAc+Y0tiXGt5ElNE5DKdx7Zoj8KPcvYbT
n0TdDCARScP5j7W3kp2/skuSi5CI+DtrBVcsGfeQe1oSSQEk5F+ql4CB6dUgZH0n8hancX8+9zkh
+j9LamT9eL6PujLC5oJQhQ6UUoq4pwPcX8g0+ZC0Z4DIs6PO51y3it3sw9sTuQpZdoJtmb+OLxZZ
9mb2Zmmm4SSWZwg9kYsNpKxkc4bLk4ViIF9pUDJE/PBo/2wnJiQpxRWJ26jc+yuxlmAZjOGyFnCK
3CsYVVBs5EZj9LODf3VwDV1XpdHKUvvDx+mSwfQUK5lr27npIRow5ALNUVg/kDjODWPYuYJmi87a
JV5Iy+nJmKg532m+6oEcvur7NS8yuOMtyOxL2QcUEnToAg8LszgWeZA+ffs33gIfV96fAbcCdG5x
1Beb8oS8UgzKnO2ztOI8mHzDlw7P6Iyyj+28zSQN5searfo00fJxgzM293KU2EOffllEpvgqSRBZ
LZXYg39vEyg+a1fZlsQ1Tcy9Cw+hzNMm+7c4HBKkQ9QpXxSWAJZOGfF9Cn+Z8OkC1RyesuQAcGE9
Q5+AqS3oht3YnhZ/qzJaQMnZLIuU3mYg1PxQ9GVbRFHp3wC5ycqgT/3PQFHm++plTC1qlyXZ9/U6
ql5inc3LoCS/i4gROw2V1IMS6WkYAp0ZcjhZp5cfYaaFrTAyLLXmJiu4tXBpR5hMYMj+x9jo4vEd
4778y34kZdrgdumvnP6IDdxeBFcw51jB5/Mzj56rbiaaR9ytpcn01atPgG1Kjsij2nDp33C60OHi
gd0g7XoxCptJo6Y8iv7MfvAuZ5hsPbhKJaZVMP1GCZ+paJZxxvsk2liD0AEl6yNXwxeaArBlkOAY
D1QghKuxpxCVjW4JOrzm+2pT6iYpK95WW4pOVykJG9UNAzddIdIC6Dfacqpoqzlz82HC2+oBgded
eUH/opEGuV3WxEawycZowpna6vox5NtbplzjI38A5wEMLMvftt6ptsAu3MgT9mdx+zVw/mh9iqzC
uVVDB5gItKjq6qV3KEn4MI4Bh0Do5y8piyub22nlZeOn9JPPgPPL3zcoJFE1zeot4fAknXQrmh6O
zjA3syQibZFs2T0KyRjz0JkR96A39BtnCYB/a1DP7pG1AVm4iOpQtQqRk+q58lFCofo5NO6xFQ1k
0l/VssMER+/Fi5Tvdwp1XpT+qObo3Y6yNEWwdXwV0W4DPzTsyHu0JsfC0r3R6Il+LoMWgjntMEt+
QE20VxTeH2u4+n+5wuhJePz2DfZ+0BDMhDuibMXtobXvWdkVzUZ8AVIeX39qeBYnbGF9ylTX6RdQ
69l64ooQ7YNt2BHQLRFTTqDp+BNmNDyCwy1E6+3aZfrIvljOZsnxNbJVltQPijRLJqOMkRRaREg+
CCt9s0lzMKGMOzxUDxbubBWtaVL4B0Hgb0ZJVXwVnY5MsvfedS5KSJVaOATXFOBdoEjVwDEJQl3K
ry7QQ6rzPTqZrM6S1BeeSRsRKXDWJDUaam3MToubPHiQal3O3t1vkoiqmd4oCsSfCk+NiKyZjwXE
sD+uQBFXN35Yq+HVPn3vUovVo3Lig1YLK31uzzdMKCiyYa/lXQacCZ1DYCnhInrCluwuhK/bEElo
01YYN2o/QSUd/uUI1m5iT0hcQMCGQtm4n3vwNNK5fw5qDCqqee+ehJn87A4uUGpSBN53LiuRwMbU
lnkIrKugtIvoUHFniwPQY/Amh0sbTo9TJfJFaN6NQE1/X12X0Yo/rLqI9RwmRpjIRYR1ro4+eNLy
W2X6msCZ24wQcy1fdacr3GA/eDjVzKHc1adSXo8AcaQHXrO/UoL+oWROVXp8nlSXD7VKRZMI7ErS
lWhwk6poS0d7fr7TK6EuZt/CeSmrrM+WDvccgNgI0Ye+tjJgyoCpBc0aonCkB+usnfoKpxkizgGj
H3fRtGYSCjo7oIPy8FE9XitVOsEP6c9YJluJW0Vsge7rF0ihYPabr2IGoEAELxjmetvw+3GF3ipt
IODbLvzKWVLdANMv9NK10PK9vr/arCXpJUcgy+71DYNjDXaRrVWLvQeBki3Ug+54s4XTu2NeMt5W
Mjso9v7fTuV6UQPMcDTb/Gr362HE4wzawg5lvShExhUvCvEXh9s6e0xepHnYH88P+IPXn2z8rGWL
YGW4rNBlvQRqLcBpvcTbsp0tV6dCN1lKvCk+5VPJSeBe+lRsJmtfOuR52rPZj7qD8o+BJYEKyvZp
+xCLAwQnZ3NJE1ToVq33Pp0hiJ5LLwTwSCdNmkaoptzWRRlD77uRZw90CMwp1bqtQYgxo62Ndx0x
w6OMKbE4QrJJPxMt4ledFhcGENBXRkJfH7Rj5m74l4u4fBQXsz4vKFRsZ9SPaFJO7hl3FXDJtS92
2S3s2Z2oAp9byEzZdvo2l0pKwQWV2AvrmnR1pc0BniatI0v3w8DlAc8KSCVtRXW4goHKRdyvP87Y
dSNJV53ZNueVtwRTBVTgzLoJnyps//rVXbYbKLgttipztCEtwXKq/EpPeJHxbXrFq5Hdp+cMCcLO
P1vmSG4IN+qcy4D+Vbn6Lv/KYP8Wy42sVnToRZ7Y9NeGmFEfjCi1Uj8jFO9IXoe5ZzlP2B5Yt7tq
/U/bF3B4feCa1ddUdXku5R2vd5xtLg5OjBsGVSonS3UOtsVScCOBHwOJzO64AEfQ6paO7oWlLfm2
n+O3pkf4MczajDA7fI+/O5hwq3lFrm6beF8kEFjqm0h0GueMAajbkStylZFbJYwifd4DvpJL0c8d
YbbZNJlFKtmyNTkp+2BnFFNSUsQA+Bimhu+HHnV59EUjMizhQaZIuRMkzADjqEgYxsYB3JZHkq8P
Wiuy8Xo2hCKRtlPbtxqJ59tcXwadtsPjScpJvg1NoGtXzEpSlHK0FGwtu3SCTkenLLZUsXiZDto9
D0rLcxl38kQiYZmrPtKB9EIk6gwofoXsK7meWHCmuDxddmvi+yTZSTtmfmCbl7taz4BhSR3ayzGa
KHIKkQKYwoK+GzFne7q9BYoG/UvMo4bPAQQfr773H2/7Gxez9kBoAC0wFoDI/I/QNCB4yYd+uLq+
Is1Q0Vg126PduQOTbub8VOUqzxmCoF87gYmi0LFV3ibMEpHBA9YX7apWFoD03iL/thMcvpJ4awSk
ihLJ2r+Two+we5I0o81OTVqC01qlPJvIHiKouwDGJHp6I+4kF2MQ+PQG6RHnclIve8A/CHjfyIbI
ydhb61Mr/UAYFvFaGxTPEkoemgnD/cM3Cw6EEdltAN4JyRPSJkgePJwS0qhleQHVW5PFDLUKd3Db
AtHXsYHPaEu4w9wPqugB2+wupOInZUZyl8FhLV8IMdKHusDMmaFzG1M0uKcvY2FrGoacYXpa/h58
zx1l0VuEkv9X0tlGfAoqxRGuVp4AOD4QYUZhYL65gq5WkEjWY2S30CzMIf9HUbou9y9J9Tinb258
/4ZlVRFf7wKDspCR9QmT4MVKuuO6+BnZjQIR7AtJQM2fbqsmqApqAVO6UdHd/RI5YGG6p1+BIXmF
kpFU8+hrguq+0w/xaPmoRkADvP/mjgboFtJSqm31gTXrlfdphLARGw4+npKcTNIQgZo/072uL6rI
/054eUZucqpbLeDLxr+Yg7envE2zWRoDQj5emreqk5+NXiJ/99Oi2ZMP0gG7sXttip4Ta2QUDH2P
EzelC2dVnULo0W5mUNlwUc6GeZsXZwEF2CdpGm5YNoOqf/MRPue30Sn/WpcXCjdluvYP2K3q2e6w
ZUAsvoCG8aEUmlWqW1Od3ul+GLPj1YSEEq8FC9y3TDsasA/tQC40A0JEh9EIwu8teFDlSGcT75bO
zZ+h04izJrTXw8XHMs+riAzSkszzItL0uxKxV90jAYxDK7ytvyoZy4fGSlhJ+7vXNVcdsLosLFWH
OQ/O4IAncaUhBtDdIQigWKg+Mf9OyZ7isRlStRgXAVPAkhyZ7NdckgM31zyv7uHLSwLhF+KX5CwP
WA9RkgPsVVj4twoPbA9iWulQdnuOgUlfNsFjFoBTXw/Z1aYfItuDGkioPI/gHQI4wMuWW0NJ8LFI
79J6BVFz1s91MaF0/giPS8wh+iC+/oxGONH0k8QYY7zSsTsSlFCZnahUedYKHrtVl618P2fLHreV
RDCiJeQD6ERj/tJh4/fabR2fM+mc7yeb2Uar1WJbgUe/veOsvUr1CkwIyOzQ9/B27PlKOAMteuo8
J8fo1ZII8k7cFiFUEDPDxx9hT0TPVjDOVHPXRIqrfkhaqGouMEFa6t01HkYvCZ6Opr0Yyc698/9Y
z+q/aJgraWqY4FUxnbMm49GWzT34nme/LtyjCVQwlrX2eXPo2aOztH5tCtp0H7GCYBJTLnQfMsQF
foDcvyaq8lsGht4vBPvQ4zdLzQg2+SGojcAV0Twxjp/AYKFuo6nBZo6rC2yPwqHjRGzakNRb1Ans
HOeUvXdsaSa48ULpxCcTeh0CoQjroEM1hJ2hJWQH9WaSlgcrjZxz+GYaL8Xoc3NaWUwYX39lGU3+
hIbBZvJhSX2Owx58qlghVMq4Cc6WxrQtVnTHV/WcfnpGxUNAfW37zFyVLdySvjUnukEckqz/ImU1
IG6OGnjDPJos41YTF0JfKbW8kfigR9ek4GH5ZLmQpC7VYFpRFD5cntyQHuPGr+Gbb4uwpQydEGBb
v13bsc1SY3Ac2iTi8Ks5hSOkflw8Ds1fb6KPy3PIGNAMpFdXjp44cqNUT0rEUAp5dOCV6jxT5MqF
dW3lWcFgmM5AQ/z6ccjj5jMbF/MSErgR0bkNzZCMb+sjLbL9uO9CZNL7VYM/gXQ80RRgLXEcLsbj
Rwlm+tPAvzzomkDsVDB8pm1u7AAqZEvm3Zj6UprPxTijC3bR/sbBusyw7nXMKxiPW3K3UERQZFBw
mJx5KRig311TyzInbWwpvmH5DMyXCXTYMJOLrPcVyBZ0p8f2DMFTHspkkGwf+55YSxipVQMZ7GMk
YPtUhVvlih1+sUfjnwH3FvGcs1/7motLDb5a0SiThOPI6X6TJRtl0cIAhxQG8N/p8eC1XV3nR2TB
g9xC4FKhn1mkY8/dU2Cz/6NZNJN8BbmO1P1E5hgMAHXc0wQczNTYvO4sDvPfHuhv8ZdxC+dePWrS
25bI8L+8PzpuJf0ScmPmtX9Xh+iGahFfFM4NnAiHm7svBMRjSKQjxAsSI2bgPG0BftxkeGLdmqxw
aVEWeJmiXgdfrE63Wcwsltx/MiKjNUtfL9rEn3ICh3kHUXawEnHMsEg9ak4G3kIMrsbKyHk25mbk
OHhd4FjI3cgBgCjK5nt47HmrLYQ9NQWMGO88dRPN7lPDpyQ0SgyTseEIiV7KpSJaC0KnXUrZmH/e
Wgvu70AYZaUHAzLwe/T5gOjatN1h7V0on7CVrzHh1XNLPZPycd8ygI0kHfS4w7feTbv3Fqcb2k2N
3K+V4fYDTwzX2/ASFYCOqJYEaKE4/PCR4aI2Hc2NLA4GxiLpDw0Y++9GlpZ2aBU5HsZzYxAG7CJF
3DPOWQPqCfJcXbAaHmsAYHA0Z63q2dfkflm+75MEErKbaX39LCrEHWYDWefBsa57wE8lVXe7Ig4w
S+W7CXnK2JX/UHn0yow6CHLZjZsmohupLs7CZ1gJQDfwpv2OPyod/pEYp4DVkyiedwKqbP2FJiQd
VicURf23evxoA497D9DzmaCBgZkFkEgfa7aWw5sbzYXeQWi2U2s/n2dJZ2svU+pimddFneTiPJZq
F3Pq2u3XXTt89oHnnySTVzf8IzXyNohCyWv+YPNE3WnbCxOIG2mijfNw2+jgTCLL3stOctmhnmRt
PTbC1kawsg+JD0pOnmv72jzwzVMgMWGMG0/wGB0ejEGjivr/EXnihhRYucuWJFqlVG0JD00gm/OS
QjPZF9iPPMXEfekaCnHqoP4OZGWYRLn0LMIHp2ZYkB/6qcYkExTlQsQu5/qggIEUwt/xP+bVftNF
HrcSmZpTpskqd9EnWIxkszCtozd/bU2kHwBq0n48gWrnXzGefXvz5bM0Fa+yDgIjGuip+YOoIty+
xy4PcqcON3GeQm2Up/xQHWdywD5CsTWPZLMSwtJRc8X/UCNJ5CT9kZh/isOTAvLKo1WPfEsYeqUj
W348SplpA09U23RlmfJVbbhdiJgCrXphXdrnh5eKap2A4Nparmuqd0xgyO98gVyyQZO0+R6YnBbC
CtB+O99L90yCA8nacO19rTQVbVAdf1/77NoByZRpBbpq3Op2gNEOm1p4HzdUfCwU+zM9WtX4yh7K
AqS/DEd1xHK9kTZn+PQ6xCAQJ/9w/zqawcqhrqD3JTLYndkoqrlGMyz6yXTeXB9rLE0sO0HzR46b
k4NGzdDGJFFhWMAUgJpF3wuhbac79trWhSK0vkKLSuGRqk6AUDmvSduRn3b1YPQD2aZQ+GOdbjZ+
PTX+NjIevtjDAjM7ftWW4DrAp26CJVzC4b+6o4T6eE1FQpnNpHs9JirjWqTof4pFfWQG33nYLiTx
L6SVaP4Vklxz8a5bXBYoS8B+65bwDNtIUl/jzheum48ZmaiBQe5bMMDiUk7HOpKYqyaqkjeHVVmr
FZXCIfr2t08fgCKG1xIbOzRw/BTCBBK6WSAWpiiNI9kQSnfuZoJG2EkJYIzFaajFfjxu9Z39JVQt
dLpSCpj+vqYJ7fmcUcLRFsJuGjefh1v2bPm2u+tBdRJfgVi4pt/cGbbLzuDCP49E/enujWOuHk0p
Z/OcoreuNV9rm6KcwJ7IbMpWHCGMNizSeMKPuDpNhWZQBHN7AUyJZ1q5sMgYs7TJzFlGdpZGYARj
ztpyvyFt054DVgGudg7r60NN6vOFZjsPA3a6V4qGYc7Bqk7jltcpQ60hObBzdkZeh1ypCgEhkob1
pj3c5irNOBZ5Gj/tYPJbQzrg5x/lW+px2Ir6Vh9yCsT/6WPxsagWeLhqkBwU03GAptNENg/9vR4C
1YnQH+K8QiULhLVRUQPY/ry4dps7kyohtlQ6s83YnulJjy3dGMc9oYTbGB8obaoqU1vpwwGjmOss
bKwYQ8tHfAH8X/1mWnGpAQBCVu2Mw4H+YPCjnkaxYE/5yAUbuLQ82XPI5SjkzJ3VFA80mogmUf9U
Vs99MmbIXY+NmijoxiP4sg0Mh7+ZrMVoC6BH4/QjLIJ614Z+AoWRCM97lCGXCfDh4V4vOPjYeEm3
kkxcBc6GM7Ys4juuTzU7ip0yoqFxw1x8U7+eFshG5jKh62H52XOFcnDSTSzKyP4TmVjI6xSM8e+n
5MKcXGFbpNZ+gSoDIBK4GMoGqehlErp1ufLwZPAULmojvqsWHwJmM570xbtekg393mexnn1cDmoY
7cifvwzQ2ZZ2J3aLAwEN7zxVr4DWuVSJXTdu22HLNzSmnF4wXeUS4XljUUcWQnMwr8zRLIexBYXa
JS1TQyAOXnag7irWCgTItt9NpRrRDA1V2JwSKAK0NJaNppAwdkY9k77q6x0umZC/MtS74T61yymM
6oQ4kOWwdA6CQSgmq8C95mbPWlxszghfEaHqb5xR7IjhO3lojafLBf8h/3MoqzZJng3/gO2tSDy6
u+aZbzrLt4aYP7aZei7q42sOEv+TdjhzVWJqmRjgdU5Gx6XQVbOcUejujhTUxxorP136AwQ4u8N8
ih5DyJIIUx+73SsR7T74dcSF7sZVW5iWElPsRzwESXGX9vUBhdQPQHLat9bQqNuLlp62DB5Z0/JG
cc7KG73gICIN+VZBzLMsEUc4/Z58ShSIkQ8CnqCPCYb3OXC15vrJKCBd3kKmlWjQ0Bgi/Yy0wdTw
0okly64NldarHRRb9xTJ2Pm0ExttP/pp32womyLeO7ANEiCorvnz7Uo+vc44UjsrKWKmGebq8kO/
+WGlASma7zgYViHgT3vzx05BvrsRuT9BlyJ/mLNenIZMjImCcX0XXWyUNjSeagIt+hKhHN/bCKjF
D2VMFzwwYsAadCsfrhzRcGbraz6OUfBz8Mc+LO15IbALRIqV36w4Fw6A1+09OIYZm4x9epkim8UF
Urp7+gGvPGEbMToB2EnxfPaEb0mrQgAA8cvI7eEux9fLnU7YLYB+3rQGBtOFCJq35g3rDuyUlh1J
iJyrQv2uheL6/Q7S8PN3NZTlf+p9f9s13C4H5c99coyfWGsfLtCx4RXwd6W8QBTwJpEHzJ3iWBq5
R3Jp5gVg7WJGnR+mxHgnjcExhIvmRnl1a2IGC7zO2sQ3I5eGVmucX7W66r6cX7biR2joG9RPrr5H
ISP3jTYDhr1Vc3AAK/OVb6BOD6MN6Tz0lAL1GqWEzMp6f+ZbYUvfXv+g1V7cieRJ7Ul4JYlEedps
UG3q23bxMu3MdyCdhfsRLH15JC5W+kBNpoBdnA0CwLXVAaLzI1u3b7s7MwKk37kFwY64IT1LQC1U
iC8YmfqfKUfGBkwhNo3oq32bGGXOP6ARRqgL+ly0/41r2/cZ2Zt43d69hrJKLdvgZLeeW5vE0+D4
kOrt0OL0ICD0N3q6+SVXRnpDSxEm9kpgeIk6CxlId+efyl36fdaRxptWud/bExiCal8FrKXcNpAg
cTdXBxxHwoofLWYaFLjy6RaGPp0rGiI3zML7gf6KryWXJYuIYodeLibj/gZyg36Quiw3Fu4CbSFT
C3aAryQFcQ0vxDvN2MhvrfCFcnDHOJiR5p7Auh4KTM+VDijqms7/J3EAjWTdd7AAG+1aMz3GD+AK
BcCF6O3ombRKUQHnIxGwLeIAxfEq7AsaYdJkALnrARBCa04XikroQATD8LI0BokFUL4ASAkLwcxs
8H3jGhaqSjAcLvWPeZpStAQ6sXuZxLM7vvmIyEuS/VOFjWKC99gA97n25B+eoinR4uJeXvatqPGV
WljIxhUvJ5osAhhGy4DqIPaeoKiY1xe94Rr9czaIVvLjuxSU+yJhavXfatZ9N361p/I9ASqJZAbx
q06HSLSs7aM8mcZ7FEFXN/i/R2/jRlZMYe0V2bXovhvH0K3oYvLITkfyAm3CFTGtE8dqBguvOzQY
9ciSuPIYzFkI1yI6ZH+OPnNbg/HNuuJmHgbkW3UtiyZ2fI15R7kDLu/CSd6dZhxDEZsAAoCTvUq3
NXIu54VYGzQolT50SLYSYNqnBdux3P1lGLjUC6fu191kwosr3G6M71hKHlvHx2ApBWaJsYMSL6Vq
UjRt6CYe08T4tcnXOE5U1hx4wBJL0V9NclIe8/+/8xEoOJkJBhv7KMrz+auUGP6xY8VsW4Ylrp9L
E4grjQpItNcxh58PnNGwKLco1b8phTBA1xT4OFRfhPiG0NYnoF1giBEnvaqKPt6QxV0ueJ2UhbXh
G0c74BUvRZljt5S9aqX4TbO+QCLsi5z6apKhXXNtzex7UtCBYJ4Ppuvs1XGY6+b24SXFQRznMofV
TY8/cM665y9jJlHcuL3zx3ny1x6iZ3RcZFNUQp6y+4bx/b7f6YhuAqxaGel9wiu8nPJHi+X1ndrU
TSWjpAXZhEYjeTmoxYPhrHYAMCQiUAkwKHDsAFHbpZ54lYZV6k6OLEIOFKzLRDqBSNDpAedLmKq8
p/Y9Izz7izoUhZIZthEeB/YyEq1E1vSW7/tO3BjRaCEAJPgkn23g+I6e7JlLInIpfNA8DKF39o2o
fKsdddgt5mJgYLFQAU4Wk9ngIKjmPcvs2duQwIwuWRytWBqELk8favZNBGkCARAu0lAtp19kpmY3
PToXqq56MtUlioWol/d8AY707DQ1cIrc78AuBNx5rM873eeT8vmYvzW8eyJWohGZ58Lqjr5pxqAP
WKxKRMJw8kEZj9xCCLtKBBBp3/hQT46Rd0mxPzQqJyswfEh+h9WbBRslGrsNhtodU5IccBxkAwql
esHsvNJju+H33pvhYVrw7btDAgI3uehlLbx9nVjFySpEWXQNMnTrRKyr0CmRIqMyPXNIXf1LXR/C
xrGxHZG4ez0GQZ6Q03rqlQEZpoa69hlEx9yXXDiTWbl5WklJK+NsdHJXyL8ifXomFhdllgJMv69w
FZd/NGZqUvppqKuF9x7gvKgrrY34dBidrDTnDI14SsGu0JRiW+OiexKGjC17uFG1Yc0eK5Wl4xzc
o6+hYgKPW7XCyHZfzzAnSvCWAZehnsDl6PgIf9XtEzm1KMXXmKaw/CChRWGb7EBsb/TNBvL5ZIHd
jWRoswq59WWfbV5Ixw9NpaSmvRP7yAIINDujr0ifzD4xF6esmLXWz+50WtvC0upYpPt3h1/MJ8hl
tdnB6VXlvRGurRU3yfIynKZrSk5Elxhokvqwj0Z2CO4hQSjVm39XFVyElyWxBIDEeJVhmXKSpo3X
BEUbUnpFf/JE2EDzj9brns7vb2UZRAW6bnPfgggl6XvFiOb10zybBijdpejQ7Sr08nOBzVXvnxm+
+ufKkbV4BhGHujaDXUPq5G3+RoRcPV1SjaZ7KcJp4HEXojIy90ZeKHH7Blw9gHbslNtVpegTftiN
rI3MmXCskex0efS9dVpblEPqotmzwK8M7Q0Syh62ohLShrqXOUqbuFCLlKKkKVXK15oG/KyjZQWo
O9Vto5ZwseywCzSdHA6KWV1ZLd9F88Rmr25PrIFA9UZqA5hcGEEAwTnsMIP1dHLp+5Gs5P1TaWuO
lFf34sCzHKrM/CnTzOI1zQvS03IzIuNrfO44StlPbucQEXII5O79YwQSj+ywI5xyMnMt5P+tXLzt
uvDIQlXr6TcBNlBjQJUYd5UUMC4f0IIs2z5i2NvjoL4j4KNrVkbb0QwQ8Z2aNZy12KUXvVZKHMn4
2oXgEWMr/11o2kE5buw0MDKWf3z1hYCCzxUFEi199LF+PLG25w+6N4KEE6ocFjdcWoYqdLgzhggc
KTo6AMLSO7tK9SrmZrLzJP7bxo9cf6/vP/rLmJswN4fGyluuoSGAZl3Cqp1q9O6j6IzfZFxCnP5v
1NxlKmuiiDSO9jVGiBBQz84F83mEvQcXUlUS/wJC5pZwQWxPqkriXAprEoMLU8kbJpmabHQVlDDs
DOpFpRe/cs0FTU6bAv/r7ckC5UPPCFLzHmOwdDVPeSarkcFrt2tAe9kd1J1TR8I3vWeeDfaqXKNC
iv8M+AtSpabEfWuJBDGu8pFoubVvzEYYvRuN+7ojvuS9Z88+01/u+LNSGQ5xvpSWq43ae9dE9M4c
CAh3PJhnubAohfxB26BH/6gqMjC+QvUN7+xuVveA6ICE0RlrmEPCcRGni+Z0SWKG6yVZdqfpXTep
Pu1zlirg5+W9EUtSRoLIXqLA4xfLlh/mG0ZagnuoOHXhRleQnkyETi1BpJNUhgEglmYuRJEXZIif
QWf8hrISbgo03VTfninZv9U0TyxeacQkpgy642hDYZ4ErgOSLcZnDiwZd762JzLcDxCU2TZjDkrI
J84PSbxamDvRavkjtmTf+mJVavb5J5OTKbHyCN7Q22oB092C4yTvyTR2qomFe0TM3/vtEot2foQl
zkCoZgIPGdUGGqozo+VwUw6DY7Tz77pjJYPUDfYZcjYMUO/MGwS1q1YruHjyIFYr4hHaID3OMxUd
TGIsRue91m6ySVeHEamiJITqPhdu66L0+Y42AvxRXTjja8mbx00Eq4w0GYNeC7MdH7izwS0n4bbb
7i9OTn3jnvA24fLCbkqlnS+2hHUVuEnn7MLhZx/+OHwRa95J0RdjB8Dg37mfiD41YSgE73Kisx/P
MEsVe5ELeAzTidX4WxAw6/bEN4BuHK0Xjrf8iCpFsPXyS1a2A5Ikp/rarrsfvd7vlXWeXRqHUQ70
rNHf/kbFuPaBvJVMwOqB/3bgjKHKaTH8J3r5xsKpd1bHGYTu567mRJk35IqNy5lJCc3f0eGNWcpb
tyMz+keNMbl40+Fzvqult0N/+ZrFRlfhcPYYqqfKna6ieyvgtK1lV5A9uIIB9JQaGX+sRqD1Pl7Z
yj4t6VIZJOEZd4s+mJsDs4hmKhKpOQKE2IDgt0xLgPwXGAoVSP6F8NQNw5MoexuMC3fcTmEs7Pkl
5nw/PVp3MsDVFDcRcWA+JnqpWj2BrOeHm/2LK56Av8GL3iXmpJPGZ7W8uLqylBOJCIqvw0GFBJ3y
ri1LITH0jWo0Ss5CK1Nh27Y3pBag1Ae+cGzOPrPJn31q7VMryIeCItIaqtRLQhcOCD4SNn8m2+o+
CHKqO48FAWiAMBCZv00raEpo40a019xqQqfhrwDfY3YMgsTdGzZL7u4A68mWGVKID3OP4mpfRVMi
0tZYaez4quWhKgTLyuwjHysS5y+LzmY2XHt1SZEWsm5uj4Xlbs7HCqHO49eCLZVjQHwhqr93S/pe
bUoDqZ6+srCk12uPsxmS+bIu65XIGDzgPP14ntYoA5Ap9D21XbVapjrp563sc6uKgVQ4rNO6Jz81
CcO7VCeoI1NWA9yqMA4o/dMmy9xliOLR0kE6gNEdhk31xejBtHy2BfQLEPYNHk360OlaYI3qn4m/
uMCdjcSGAO8FogwIGBGkrmB3qfsn2OrC11cbm74PPF4YbWPVqTkcyHdlC5e7fijrEOEbt41h1GLA
6Kz33A/EzBaqGUQsCvdhpS5Z6R14P3nhnD1CnrH0Zby/9b80QShamN/njPPYW2k7lL4HXJlmkp0H
5t9cjIgTGB4m1wN6x4jFRBCKscvsgOucAG9pP0c5/zZnicWf7MdnQGWmVMgo51ldBfxdayW4MIqd
WKpk+Vx4QBkhC5P0yn0dr00nkZp1tWpUWm6UCyh93xerPWuUwX9bpZ8iEaGLNHG18faBbEMdk5sS
vOZ+U8sxRubhimpl6vytADYCkW5sy71bUnQ/GdtSUJhm4GHHwJjsmA0yPXOkv+WZ2PDiYcc3cX4t
yz9OfzATWseN4zCr4kteB3gIoyycjNlQKx2i4f28WszC6gLcyfuMkkThOgTOQVzpxWdnZ+NnUVFv
OpkzTPOfQTL/LR7XlzP3NvVYc+XN8tJNXkPzw5bcOZj5Qtw3+TL+2aE1pKjosMARLQPqq3YlykIS
ecDGE2AqG/Ppen5P/B7V5YJIGKo5MXbdDNirBTEQcjOT/kydEnx5c4eaF7y8bPqaPMFH8jCOZz4f
0YAGmKH5fzH09+bgGB8mlVck1CY/4OiLvgTXN5jwWt428Sbph3nIu2KzpksXSVlXxOHZLQBEcS5L
SqhJK9dxGP9121gZhP84N+RJwcDZ5F1UH2O27HirnxvRcjLlYIaysJOkMZVJRkiJsg/6lObXFzF1
R/iN8X01QvXCKq5ZkYYiGYiWeq8Wpcew81cMMjTrhjHWM4u5xiPiJOCrQa5pcyTsPKPbe4WewLLq
+Paf6KpmVQqwdPXZON2RUW9mjX5x3OFYvMMNGqj21qtzgb1CSrdPC7yLtGIhP/JL//WZcVzH2MOK
CFoXYAhXB5dd+CLjHDbTKR8ENw1VzCDQYpCIrl1+YIF5MUGJh5vvPzB+3lW5e4bPwctIA8uuBIDd
KYXb95q1KGZbgTXfJWaLy795zco6JnKTP1xBaOfrTWXeNCkfywcrYShr9mlWbhe4aRxhi0MXhIwt
IINDY7qmo7nNqaejyAOUluFYLphzSsEFAbv4DclJsgayzUogdV+uJQdF+wLmdxa1hv/yuCm8jgeG
uPXh5Wj9q857lxoAPu3QNVYAHtkXu6h0JxirzA3UvuElf7frqPHg9GCnn9V1BRs9/qjeOPD5td3d
3LvYhQ2DSp2jLFWQ86opYrp7PmPEjXAPp/zqtuIuDtH8fkZF2h9L3Hv/4jUF1akCaTfMiNJLkwNf
VUECi1DR1aanQPABo3HlQxE+PQwjqXTWrkth5eRoW2cwl8hkjdu1Vkip5RcPArXY0eyNyd1HYtr8
6duX2ZDDk8x58XqHLrxRqA8wZZqI2aw5ZoZkJWvhI6Y5zfwy0bAOZCow5+mw0LEhBEh2C5P8aZJf
RyDHGzMD9K3NR2Ep+1BcFY4mCxkKehjdE2n41E9R3KTsKJUrLSF3L/Se/onYYoA0QMrMxmE/w0jT
XV9A07JLz9YQ4OMW71uTHnXpFhPcHyzr47w72lpvVednK7ycU/q+IlP77rowctkx1mFHEfb+0vwP
jfe/t+FBbpQBt9f3+mPfS3EvAbjxcH3rmaWm6Ni+lSTH64w75utQMmh/4hFWGzhoGcndf869cupC
ePTBuLyYuryhleOxgYGoS4a4IqvXLSwcK2Y1NCbFYB5WLuCOzJUegUsg+H2K3qHZU/mvTxwcv4Q2
DBCK7kV+zM4c6NyjW93U6BHbZyL+itlmBxSVWQc6haci049oIiKHGixb8WnvETmZZovJm+SDVpyY
+OOljbWyCd/q+0zsP8aiIPNmWaYWYXRP+H7QtEioZ3MXrr/e9uqI5YoGtxeV7zaETymnEpGM+0sk
ZyohnfP5rxrCvuXI2tSNd2Ka2+7eEAAdMLLYvFdiplSMwTaaE6aMCwaj070/029OfThd9L1vEwKi
9bynJUWdOgW8TBOWt6OMHc0r2NWfK4OwruqdjVZySEXh5rdKcutJgoKvNTMaiNTk6RQE3L7a7Obx
DnTmAQP7gpuuZfS+niXVcCOjzlz4zt8FY5mKtTqI/kNIn83JxQzV9EUIj4eW0K+KCVxjVHw1b399
EqHSntZKe7xw2d8TVoGDj9yOuUfZTDPcPXQE2wQ/fOn+DnaKBbETT5QU/mwVJOxhlr2aJBzRtq9K
SVgmmKzC6OB2N6epkPxc8DcUHCQetduw3SNtD0I9sClQesrl/WkflFzZLFdeUn4PTHBRas/k0LP/
EDMyaisC2q3vNG1UTaYnK0JV1wD4lv7OakCHViBD3dFL7viux1D4dGWbRaMYnL0zptM/gK/n9Gqc
UM5bz4z9QEhUFmEzGDEXxjCR3EC7m31BSgPwQsuw1krvqCfTAo+G1ZFHxIu1WWCf7jyvtwzRr+1p
Rm3UY5EQcDBCB6AfkifkcqsIBaZxJ2mAQxcJIKatfO4hI9vRd0zGPnEnfOKrsKA5rpt/KYVsdI33
w7wTaoDKdmzyvu1KdfXM+/SnBHfxzcLE3R9U7X2NY2H2fW6+N9A9oUFNQYgFhzwqJobZmidpuo8C
cjiZXAd2UUhyLXSS7eR+d8aH8DQ9irIQWARrl6Oh4mkqDHLKIb4H+b0Qox90upItP+qkIsG+UuSm
h4JEaKWCjzC8oz6NNbNvzqfvrYw67jhHgiyULbuOL+aPNBFYLYlLIMJXjWi0bPAhz4ymGDc1DAs2
XSnsIW4WRD1ejgsz2yEhuiTyOajiNoQRE/tT/gfvhl502maxw8x6+oMZ+qTF5Vhtg4nB6EEjahaS
R2dlvxYkp1yfOcxgVswHrNPHX0ykXcRPozsN3z2dZQ4XNwZS3REYd8OIg31JglCfcmG22SX4Q50z
xzWAKW++ebQzfY8FId2CxzNw8zONl5nsGAWRfg9v8pkXjCr9m3jVA0PdzgH145BsNOhLAm/MT+mk
OY+BmFVQfPs7GSafPrccYIlTYe87IsfggHFthSrWKDX6uLmxvQBdNrTJIP5/J7YHDffFj2SW2XDS
JwAvgszZ8sRSXNSyTDy2Rn0dA5mV3rqUa+xGNCelRC9WWtDjQ8J1LSYlIbSaxvRkLblrXrgd+fE2
HxKEASQVJCOEJMtxQvLKD34j5kJTxbhAzHXy7k8BftmwrodoZyPz0AUN9qlfPEt861fet33U66To
ZZTtR/kSkBHOT51cy+/1m2mOUetk3LeYxXsNxYsfah2f/p4tyMkFphenzmuiqj76D4fuRFTgCC+f
LqntKH7drq2RrkZHoG8Fa7V1ZLywYhCqQJmZuI53Wc8AVIaBsW+NN6Wz4UVq/qBytBoxesUvUpIH
zjEwlHBc269UzRtGd0W05uqeT2tOtYli1iU90gfRUGCIaCZhfZjx1NhfdKWieBUNBjdnqJbcQDCa
FAC16G9gPk7gFKU/D2NQGBCnGNR9MZ2igYpSpV3dhtMRmvDK7hXXkSNAiT2IQ//8lSqLRP9nmHgD
Nfov5oRLzk3tXsNQkO1XOd+lLs/NBuaMPJIPSnqgQAJF/8SSNq89cGNYN1pXaytuD9fmYriJCGiO
sCNQL5727KOjigWjaTWMRMPbvAiKOUvAZEKwLPKvu1QxXGECMnCs87O/496uFy1i/f7MOO4KI7DY
Uh+Ka1nYFuWqwonXnoJeZQS2G/Y5G/mImfMHo8cYjbOMXlf4CuHFQ5U3+21buYpSLXAEMZ1ncEGm
O3YPkyCa+nHCB/+ZugqQfui6sU+DvO1PhyM2YHP50olqBWcF9i/3p7pjzTGCSF9rgnrlQOx/dGvh
bwtEwR9wsuWse5hmRc566KKugotdT15CvmBeS57N8UAV+ZNnEZdjogN/MX7LXOgwdbD6kdKIDBZT
lHmNoptKZFfSeTssXLYB+wi7edViXjf3l8gmgjZyUFcNLKtNcz7IMz8QP2s5uY8HPCg0Qjra+TH/
hEcLWBG7mnYu5kJJTtq2dRFRqp1HMMCtudKaoFLnCgL9SDimwEV0W2vgMS1aeuuMMSxa1+C4Cuw1
6LTyRj9YlJgVaODnsZQ9cyktc4MRYxG06NYW96v1Dwhp82Zs6MoB5DpBbbuUOsrTGkB9cn2HlL7N
qxPfrWg7K4XO3j2gyZKm1sLWBThuvQYWNGWhWVJZ+5kw+dJkjDsgoqaLW10Z1xm7OQdLdY6r91Rh
popNUDfVSEnN9oYCKeZwhEKeSSqijVmoF6J0/TxOM6nCyqqlc/h8/8pKND3vIGY6txs4oyfpunOe
0QUGS1rAVLvkGj8l08aAka5xnOcFHnxwu694L5FRzcQHtqHL1RiX9SXyRZeeNvHZLvj+1pSGDvva
0fmr+lxEsGcvmZ1VeZYlGI7394JeIkCHzkIcv0GdVWln9gZYs4b2nm3VtrEiCNKND5qIHXd3q6x2
1a96v5Jojm/afO/n3vcGuit3U6xVosdibdRPHcOQ35aeShALAsABA3Fp6InfkOyfmRGYU47zyl13
9VmSl7AdcmWQdh1oZJV7CclTeS3y271IspKj1hpN+IQFrv6Yum/zVd1QLNUvsrDzSKUTUX1eGwW5
TBRM8HjT9zRvQmdODdSAebjmh/463DqfuAx4tMsYboWOIVzpfY55id0cLGQPFMQs471CTWPws33p
Xfu6tgR7EA1XmFDR0lz8p7cql/hQK4nDZhxwhL3wu4yyJb03JNnjINGoSL6ZhTAKzkpwIgZP8fo1
DaGF0eb++EI2qvZo00LlYhbp4pCTUMe7APmczwSiO7wYjCd215kep/5YLrQzKLC4o+LxBTHKeEJO
4wUks/NBJmMOgS0vTtrjZ/22ZkoDijEY+g75UT4Q3gqDi6iBatf6XCwsmaaSMyIBWZ0esivlhHRe
xGLQ8bhVT0jsgJ8dnxGeXX3UDRFSWMadqJIlscFiWeIrYoVrn96CzFbETVWRCU417spfao6GvFSw
KywJcalJgqzJJLvbizT6pPJ381bs9eYigH3UFY0Ntj+89pR/rMpAoEzE1f5LYtdzw4FPwVrIui2r
i0UXOZmHjCe9HjJKbtemQeJBreAOkHTTUCJwuqXOzXJZBp2cPwX00a6Smv53rw+fBNJo0uOIg8Df
U9QgqMTmhUtTBi25ho9DAR84+Q/Ed9XN7uSMny8J33ZuL8sBbGeUv+i/KpytI2PdbgRPwOGyqlFe
Mw8bgyvUgkmvoGyx3kjtU1fzLAPJ2qbtz+I90imOlqbrXow+QYILWCafTbbb3xnp7Nz+caS8Grd7
jgNF6KO1iARbDYxI4O6TNi2wSsFs594WSEWc9oRwT+TLXvCIYn6kkUUddxMzkrSsVd7lMEM6dfam
thbHuYzAsMBn4TQFbYEo/lW0JTlIKqXuOeKsEqClhHaHDlUcrH+D2xDIhwTPBTE9cY8Pn8yJ4H7v
rfyS44owOmpIjf69ygoKxH6gfqhkubFBbbTyipv7a2YuSw9gn0NYRtitfAA/bIUTgqc0fTPrMkQc
sRLtrCPMDqfXKSEPUBK81fB9Ai3VLdUiIyyDQ/PKQWMlWOdR4DbcxcSizE08/MJ+cNLPetqKRU0Y
/OMAV7wJlXPw5Mr3X/EFbqFrUSL/vjT+BiADnbh9G9mDVaEi8aPQxJ1b2XoULDr2wEOo7hk/OuAP
8Egv0UwVdXu3y21XuDq9Bum+GdbcJLB2DZ+KLMaDWfAB2QAqnKAHRXMiPkFZYCxTR96FZaiLMP+C
FH6gty0TMyvrp2dYQUWMVSZO2cNoONfzdtquoREE69f2W5NB/oTwoZMT2vDYFgpJspYGfwuY6HxO
kX2OWJT2oV/1u6L670Eh/lGos+oqX8M7FN5G58jCXyXVtHOJnQBMPfFbuv7nHfwfRRmV93DTti76
NaXD4zfRZB0GsO4p3w2/YLCv2nDD5NJiqQIbWrJBS0ECmWZuMj5zwy8ZiK8DOyzRrL4dquW0UqWV
ntX3BrqiBQydQ/pWxv75/zDtGPvd6Bw24rTpcMljoekC9oAN33CqrRuKwg0l42OHnytRvFAArws/
mEzzS+Uj11isMmmtfpYsT94KdO88j2Jq1ZGq2O0eeaeF22W6lCl6jejSxUqgfRhReIrw3XKf85oD
uRbe8qtVbHUMNTn6n/YmM7T8MOWY5TWp9EFrKeLnVLWZBhchoshP1rIq3c578myFxBsVlT17ZzLb
c9l9OY8l4x953qVKRYm0ReO4rdHkWCgdO2s3Ow0VOeJ2EWiXSA+Qc7CD3aZVvzh5+iR41abHD03I
W1zXG1c6WARiJwnFO1HZO0fafuL/kQlGXDzKQyyXxOts72uMwm1U9PKjb7Scwnz7Z3OHBgMQfwJZ
WSUqv3UYobJFGus4zpnL7MFPCiVbY1vB5oBHaCJirg9nl95y6/OPb4JRUEFSkjF/eink/khh4twu
AFSLWy53czN2y/X6+dbKlzH1lZTyxORADyP9Yk9jd38Pt0+ywA0fy6RtoVLIUzMWn45rRQ8+yWaN
O7H2+tJ8GdNiduO4PnG0O/pA1Szl3HVZ8frlvKMPE6G/4aPNZkh+8AiWHz2rkNXtWvDwWjbVFZBv
G468YXTCMTBMyT84MJWzKisABulVr+6hJn2hoKZHS4eohKr5BgJp/BQRQiQklT4U3xfvvazjN4bx
AuFQh1CmcXYFgys6sEvggA4FgGDHdaxDzYE6cg1gZmID8wXtBcKJLXBCpGavCELXUoSvYGwTTwkp
gMeDSLvD+28sC0Rp68PxMdA+iBriNXfTpFiOdINkaImVStVOsg/FaR04gOGVNAkOrcJz5AAUNlPJ
GlRW3EUy1zMY5RQF1x8hWuI942b0yquG8e4nrmsDwW598MrHDnO9b9zZ713alRvlcUyGJfRaQ6GN
pmgbRdYilawMRwKl/ku1v/vb6HBfRPdCtjAM1gE0gVSYvFPmviqmP8etNjAdBYwxNFpy6YD5czPt
iAeHERhyc2PqJa0u+eWFI0S3r0H2bvfgl5UTJ5z0/20y0lu8DDpDBSAoip5aJkCkTZ6IzNozAeqF
TOFGwpeclUWPKGWDFKS9tx+9Ok5t+YMzK+Gefi80dRWJt8Rcgf2a2pHrE/fvx/2rng/cRWd16Ayg
MFXHwvJui7+DA+eQ/RJHYs9ztvong43J+/Q0E2v/8nBu1cBzeprDT2zEANeoaKA8IuqTS+5FlBPz
CUOSNlHs7InHE5NbgDDLbNIQUklftmsCfUEInCH1phAonbHuW/lpqxHIxjFoh55CnsdpEJ4i5EvC
i8Dc+6AkZd/NJZQsDM0Z5bvKHxAdcB6+gjdU6P9/Bp3kFNa5GemNwg702c1LNEX10xUH5+iXfE4q
7GgG4kfTBI2KJBcxe3y1PZLRYUdgREYS2Ll83eN1Lsqg+srQsLaKI8NUUZTh65V+okdqYVUwJVNG
d8wU9Pj+3SbCSsy/etArhzDg3P7Z4Q7LR/ppBc29QB5qKZnhjcyfeHtGlLi3/QmAsx1CU7S9SJmZ
40ohKs7fLku4Xy69dgMfKxV8Wy3AFdEmDqKZiojiP/hAXrlKPEwsXcNBW4I0h/tV5yzQnCIhvCI8
+qv8OX9FQ/fmKVx02TbRRSsiDyRsfWqqR21de9kDM/4FelxxGII8cuTd35kVfEZy+oX1nMx30Md/
JdV+xd5Ex2L/HHmFDs9Il1EcQPoRqnPqJsHMAIAX5GzPkLooN1SjqGneK5vPTp+SmI2CXyeDFdES
SqufPJN2M6jqzXhbRKyZcJXA1g+a7EeDZ6tFi3zT2u9Qg6jERx7BZco8e86hslZ/YIn1KT/ocQ3/
84gPORvjueU5jdh1jQ2LX97D3dnYjO0G9mcN1ijcBsSiiJOIQJVpYZl1pB15weNrlSTlkT0QT0Pv
JJHLSRA0mMq7paIRzLO493/uUVGKC1H5Vgv0fpLTyNVDv2u81iC1DiaIoL8qx5+XQ+kmJxXj6oRj
bA1olx7DhQikMo/GKksAmeaxTHYW5o9ZJylebkuLIvhnkwXEhfHNfVjtEPjMaZr/Zk0v9lFe2O6Q
RvKmoiJh7syPMQmMchT/TU4BSENJq0a6m5HBv5YkaAqpWUdF7YQuDNefqC+hO2Vhz0Xk6aVio4SC
5a317JvrWm2BoTsEMhzDf5G4UCTINjA90Mtsf22yPvMQC3UVVtqo/eg7v/ZCS/LghPCS/u5VQm15
kXA6GTCVGuSxaHAgVbdEivIdWrm19QTvHi5aCxhXXsxyi1YbR4bi3qFkgt4D43HwrJK9P88hugDS
evlt9UXThltIMXZSnZsU0KdkfBWJ3bfCK2wYMJp3Dvwm2cWq4NAjk0Bf2qWQ8KLXuftld4CgDc2L
9QJmYY6cTPl2Jvdk6AtvPd01DqLwdI8zgcdMllTJAR7mH+YBXmndDQAlnYFLaQmw+4wH6VXHcyj1
fCJEtEjaApDm0ElO9bOM/PV95kSzI59bN1/HXqWOhj0q6ukLim+uJ5QCKFtq91lz5BGnrXWx277i
svftKSOD7PoKKGigUTabV4aqhXgaIn6+2d45pizR5waLvYKDyswSZl35o1SgqJV8grAHzHcbiEC8
Narr7BI+f3pN+j2kqaGBuBUSCHZeoIlmtvYoz75iM7muCxvnzYxbsAFszw4torsRLBvR0/W+CCAv
jiunEeWhYB0VC81wOg+hSRidD3NJzBrOvSB3klS4qM4dzlkQqtNTVifXq8/zRnSQH3SVmztjE0dD
/ZS2ROqG5ATsSFS/CkOSMulgs8L/06+kT0262V8RDYVwGM+1bZ3JcQ2LjPHw6Bc/kZ4FZVT4L+wL
h6dPXeKCNrrt9HYaeRS3OoaD6axZHQ6u4PlGfiyPZPZ2oSpOYewq6Mwy5J7uRb4E/frtoZJJM+vP
WHgvjrweu31wn5beLpXFfxq+oA/GbcrZxC0xMPmkY3zihbvmgZ5/gtmgAY/piFkkEmVqWmjpVxz1
j/rTdeQTWB+bQPbfXLA4AmOp6mggcPYfLeWNtvmaFisrgioVmZs7uMyDMXjq8qWYSxf/AO25P6XX
PbpboNjqmyqX6Tpho6PmAUB5lOkXLp54fNo6Q2Pqm+JPRuZhCIS1IRWicMNji2bRzkT1aLRNJF0C
3tTxbLDfViyw+C1RNdmJt9x6sHgGLB5U6RIjSSx7/Yir/AuATQo6N5mU84aFZAXpjyB4NMDf4QYq
gAtm16fv2T1VS3K29mdjKJ4DvHv8OO0oVvafZiyjfTv9B1BgzBeAGBxFXmWK05X+0XyTiKnyogks
Gxed2DluHOyKQeSyIC3CO2uvcl3YCmqHAnl+NoLmYa1h3mVAsLQKb0gb42YnPzaGp9DtLRhOCW/Y
H7UeLAuRYa7ECgOIGWhySXrF9t+N8fQoD7uCQiFUbGuuZ6UB5ttcpU5EKVV81iHBzKq4H2sQfe02
ZKG/Hv6B38sCLsLGu+ufdcrAmXp3kd8uNVFUSdhZEHjdYKSjmDnmJ+cHV+VLywkc/dt16YTtMYY1
3lvyUww7dl6nle2NPg9QzSh8fDB+jP/s2WwomayesJwJtBxz3e5sEu/mv1qCPzJl3SC1ZTO0odiY
pm9pU/3idM/46/yJ2I6QOvL1MHqMdglVyNkzOiJ7zf133qqEXQU93ybNgTeSalNxfiCaRsH2Y0Dm
RrbOzZm40S6hEukfFzM3JM9t2nOD4Fx+ZqVoH1ZSJS6hk6UIuiW7//jGVtc2Y03u3EegW3pCWCzw
hZdo6A+dGMM/EtXEYG7TiZh1AqZXDkjiQkbjw+m/qQeKNX3+msAZN6XPsxlfqQsnQwsNq4i02w/E
qzkpRsRk7zukhRnVGovx2e6JnKOIHERniaPTDe1SoS7BY5Qalk2S1PnSGzGhG6NQF8VgIIpH6+In
7jvf4q2zI65L/Un7ciU31G4Ltba1P+Poj0ZL94qcNTGbe/ao8FWlVdY/8+5TWnmH2zPmugotm0Un
Jym+R/QSc3+dwBPiVcjjW2DS4U5Mhz9lolBmHpO1uMnLOBPjxe/O1eQdlhIUEdDsGE9PlQN5Oz6I
l3LHCooM5L1T0LTRWaNUMeepLhM/bpn10Noz1NIGWlweSg8tnO0JChDR6oU04tVEM7OvEa0aUdxp
r+6+dakEKAebcCxwwgoyj9BXHF0/uwpzMhIH6zNt97AEdzCzFEogHWY5y4CP3hzStEXare+OFlJA
Kgf0WhpczUz/sWQ4XLhDBSvxvilG+V4n0w+nrh2goLjBOGaMv+sGWCG14MMXO+19gCMdEsQCwzQP
wAK3I9QgPmIU0s4+ZnPSudFkm+5G2VZbtk/Wopfb4akaUTTmtqCi/p6qiiIz0jVifI9GOTJVIUcJ
yoi5dtzCwORyk3fP47DFauKH7yCYf8HoOFxEa3bM+kmEWEt7Wbi0W23tdaywKDkoUtFs8481pQOD
ippEatnuQP5FBcBm3uA2COpYLYkvIr6Jb6ROJIUbplsGANCpWjkfkbbwedNFlYfCd/jCtLfz6m/k
alEcVIya/VEL91o0SDk1IiHbncUJSOekml7eTCBPveZny0EBgYtGv/GWULG8H1JSS4S+pJy0I8Qp
zih6UudEwJZsTCtWsJBXbPcNxL5rG4kDbeJ8BYG6YUXjxOPRVqIGbiVHL0qjVj6H7pCdlkI4L0df
gzH4uOSPGbJGw0Y6Ta1CC7pTG0CZO/vso7v9NfQWQwW14f9gi+ZNj0Sb6dDVsmtx4zWfnUsioZfQ
Wthqqk3FKUuPQdFcN6NGetBmu6GgiwGeXFq+mHXg+BtcdxW1Mch6vGj9DPEl4/f2R1dm1FhpZ7Ol
XPBDkeu35iCro9azeKDNuRyxFtAj5gBCp2xgEcdGBcPpM1mObAM/v213OmbxldRkPpLJG8rI9q6b
B4A3L0Juht8TbImZ9OaAMmV4O6Oe6SBCHTnEZpe7Tp13dZfErCp5ywnD3nJabgCvu3k8P1FVTvE/
R83VFlyxkdOjcBW3LXWcvfSumNQzU0a0g/CxQw9zAaqL4ivzWsW6Oy5cMQV+8rf/bAQ26AWsizhZ
X5vpm739woAMCxuWzY5qMCdA9zxQJzu2jjFaABtLKAmRpMghZkOdJdRVTB5wWSFqeOoF/HYFnZob
7kHXysqJuqFj8Oj72/if4vWADXloRRjniQIkfN8lJQaSSqBrRaQzWinSbPOZHLj87nm0Ae6jwfsh
RLnYmTYGg4eX7BcuDEI1Cts+9fIYpOiTeClnpNbbiD0yh99y6Be5NZtBfCckXn0CNuCrAvIcXDin
yojUS5ndDCGUDlKpBp1KID68Zt3fvM39luIwWvUTGy14eo0ibEyeyQcChtMXZitEXd1dbhn8EIwK
aRuLdehO4RDeYVY+Na1smCJsA5090zGBsPpwRBpY72H8sKpmGqVW62pBuFAobR2Seyu0ibh/na9X
mnwvKIXOUpEWMt3tYd2iUVMCJaQUxuj2tMyF0DI8KDWnnPck30QKJqFPQNX0su976QjOAVjCcdwQ
JO80dY8YJs1MX4FVi6KdyIHRRnVGO3GgRxl+EtJ9AX8v3+dFH5TWtDbGsqFHLdBQeCmN3cIkiEnQ
dSOYaXRRM7PuiXe92IZSk5naoHfdbaQ2h0TTkAl/DDtc7IiFKKBGFXRg5B0LDJW1zvKQeWAZXi3n
ZjqufHeyIJM+WpG+0uKK72lHZll58noDrKc6JArd3NpVT2KY0TJEVugTPBKPnQmQkwtLg3QXmCXC
f31D5OsMq3SaDGvvk3pC4IwMKLLkbGVPkM00R3vYL4RQGJweB+waWn0M+r1sjZuPjKFR3rVNAjTy
ADWxCAbVWTkwt/fbTtoTZNHaMMRl68HgcGKtiEjIEaePc5+llMxHOOEuPdFSFdwuOOYJJ71YgKjY
W9Reyt75A8SXEywSCqxgFvSzzQ1N5v84CGCXcn2Bw8BkHKh+r55Ev1r8wza51wDBmQfyNHbZeCUH
wCPvfqV6KqTPmyFf63bfziiNAnMEHY2tCokIgBNIuPNH2kmW0D8EhRUV9j+t8NwK8uwR0PBcQCIf
0xXYwWTn0Bz7gVtxEELMgMSEEZ4AKBhqmGh+32NZCkgFbK3zgA+VVsHPcxEQ0QUtIJNQV6kjx1tM
WF1q0d+G4/7dagSUE7lH7p3bO/n7LA91rAcL1g9J5qYZU59CiZ9NCbfHoXPk1/fEYvrKKETFungp
T/x9JcZBqe9g5KeCHu1btVtGarE+g22l7ZfAescEwdGJtUp5pulAF3bD/b0/DmGBX8M4r0QXXX9E
x3uxQBtmGCLhYL+faTGOmY+C6JIZnRNRGV29Siv5odlaWS5Im/QUeGURpAvsoCne2WwAvt12Mjvd
1zHqHLs9YZjXupPvh8tH6kQCwcE1F1utw2/fZNbMMiM2P8N8apCgopnfTW7bKBBlBa6T91SqWR0k
Q5NT0+3fVN00Z/hNY1FjObObuCm3hJLPMKr5m4nB458GTWmfcAVXJVBP6wpd7slnIIugskYYz7xA
iI3HvfIzols6Wg9YriOQA0jdMBntxxiqzNYuQs2Rb58gOtL0e4CLSBrxm6SkRCJZ5UMk3Ky2kWph
Me2UkHlGd0ocWZ5VRs4pKIZ7LsRo9KJaTXeUPgXXmCLXkVnLRowy/LqFLZaIMspAH5AH17DwkUVg
l8RNiw/6dXu5+VuODItaaDp9Al9bdfn/iPcjTFU60bSTDhDX8A5y56AWhCrBzCYm3NXsv9G4aIB9
4N8EHs3xQOr8BJYWO4lB2bax1UtVtE/aZBRnEm2ke+y4TrQL6z1b35OD7yJxNUN1KI5IwQBn5VVN
zGbymWeZ0qjH4nApbbgQp0DqdaDleMWBndqfC2xPZGk0yM4P1t75zIQiPA0uiQy6iPw6HkDjGSCn
om4IumAMnib5ksfsQDy3HeWAlChfOIYCpvIWhRjBcRyycl+9vDFeXKdBBv+IPCesn4jrUFX0ES49
5A6ZF2sJozLjVUSEKMm8o1ghxxolzhFD55s0dAkKnpEiGyxMK5JP7SkjM4ycd0AxKq5O998ATwTx
9xv/i6bW6w2xscYwv91Ux/RHAZbT1hpFzC8ngtZDhlzNs4St4Zv2NjtBp2kwkuFh5bBa6VDeLBJz
Pzfha00QD/vRWre0zCKHsw8PZwaJWO5dolmIbogIixGS8zYSZQIK4qnw8FxkuoP4M941my26vLjD
HKVd9tUkmC6i8XmrqOp6IIviFb94YCAuHC0lx0fPlFUwpUDfxZgifcUms/audlgas0YFbZ1urspe
UxZK/aLaHfTzVO6VHKCEnmCvvsY7oJrnhCidQwUz86lKocRvDXbXV66vnhcpdf7wLYIpzGBiFJrN
Xmszb3735ydXNc62SupEaraEKf9d6wR+PI7hSQJstMMk5UCin1hgb1wuCXW44B1mC70Ec0gGVTEa
91Vl3sPM5nu8HEmxJQdY6//qx0R4064jei8G+lv+77nqQ6bSDTkHPEi1FOfDBfcSMlHSekQDs5vB
sBulDOuI2dpdXjtB1McOCte9lH/zUg9vzi7udGr+EbFrQG7ekGznkl0skdw8Grf8qBDXeAsglO6X
DzZwYCuvNyMMTryxf+2HrtKvcIDULegKeNc2jRN19u41f39GpUtM0CD055oNlGOc4e+PcZ2ySDN6
Sx7lCP7GCrWErQWtuqq04PQREkNaDym7SkMU9cLJnLBL4mR/LhR5gwr80sO/8HMwtzH34ugnXulX
gwRlKxHwgRgRUpFSLcX4U9jxXTDhFb3qUusZA0D/dBv+sJ2/i7ZEoRD9oWzuwKHFDw/kpZpLgCrR
kzN94DfzfcbUJWkir4vcfANOS+GjWZ0jtn8Dt1nh9kvKj67QABGz8RXuSaTwC+/GTgIbm0jGbJN7
W4/C0Febe2sDAguP2veQTK9LaGIVCHq5XK74LIZYESLcP5w6HHX2vN3bvLZWNUSav1ZVaNJtAIW9
ZeGlxR16Q2OKWhQBluNIRn76rMqkNxAvKAbFQjFTfOTNHty0t6c/IeOKO3pZzeqbMEDO+41ozbDc
1CtL0FZbDGFeNNl4KNf/Pz4JZidzKEZ3lXaM+oFW6LharSyfpVVtTTSmz3hAN45LGFkdpZwtbVSd
EbYk0mdy5KRqpCe6AlmITUM9XbrgudS/Q2efOWRu4u2bIZZ+Xtz9qGpnm6Z2TGjUEIVybmocKpGs
QWPWMKDlWfyYVupCngWw+unIxm16LUwQtNKGyiTUqI/BHx4Y0Iqf4v2OCWmcfIZUck8ubCQF6wkt
91F5hV5NSf5RCNKMi9L2OrYWXZDbcFgeGZqwbdOMHfKKNkJBnSqLcyyE8XMpdXXaBdzC2BoIZZWq
9QkAZohdVZk98b5i3S41mJAJh+I5MhPyoOXITvuFRqp87PzhL29gslCvict/fmsn6um7EjNpLSg2
O+TMJEoEQ0IoyquBu7AtaDTTGeuLkJosrY/nvhV0NbrIlL+Fzu4EA5fg6AcTD5WgI9kCBi1YII1S
sL+uibIsMrvtNQCBp4SzKpuN4QLCisQkUbAV/zKZPTAoFuE0guhTKOb/+CbYq56mAdcPfyMBusux
v652zFJFV64uSymPugVYP+FyH8aclNVjd8VmtTjLfBdo1f5S2RCgQhL+nu01oQrIYFp1o5JT3g5e
p5AEcpyNAsw3jIUG8yc5S9huGzUiaD9fAqIxTPpJCYPi7+oDo0T4A1HWliJSIgwaFSaxLQSjqdrB
BkOWIHS7ABNbKIHixb66NcQYFgI3KEGaTkxgHbQmC6cSTbu/EvpPyDxYt603QvJ+DSZ7Gx7XArO0
GroxX/sf1v3LWyTyQY6KySzbAjs7wsl7q4YJFgmZRmDjiTeGnPQPE5pppP0x4xmVdv95qCKcI5Hi
CVmlkUcSDvDDAwrgnypK0kZwjVbZOgEG9xYGO+T9k9zLyKZ0uJ/WaKU5ENwPLMqhPzfRmuFHtiP7
PneZk7By45L1Se9VR4READzSdqmZP7u3DGQJn5X9MJ7Y4vwe1ZkDV4hV8omKDtk8tF2AZ1iRDK2Q
Z+Pffwh0YSn470XusHP6ljlxvw2HP6pdNiK8S6NRvVcWK2C290b05itYnoEJqnb/h8vHFF8xSGvA
Lza4ZTD6mQlMlBY0nqu3uiHQe0fFOpKwXa8EtG4Y6Z6Sd+MULMCndsZT94usfXwQObl8FQYmrY03
9b/faa6OGr0MyQcwvUrh9ZT0pAeSzGhLWOEcCZNSY2XzReDblKs3oODjc5WbhlO2Zykz21leOJ45
kLsrr1JUA37oCGDtYbAqIdbtJux2Kz5yCGgE7MNc9bjPtstNaDGZlfTHGimHNr+divylFN7m0EzI
2LBvcBb6wQ6lG2wVgPnYOuf6gq9jMgEb5bzHjW1opr2i5Wxnqfg0AyojLmHS+vQSMAwqgSU0+kaa
922KDgHdtmx7pGMC5DZsWSTD+bJFLQ/Kb8po4Er9H32KIMjIo3uSx9+cySERZ9WcnKMwP8tU3iIH
CrdZneidOJxDj2Uz68VZ3m9Kuviynrvt4IN4AF4jcqNHjDXtI9mmUT4NVsYqpTG+jKbMs3qm/pRT
icF14u04zxLEbo7U/cGymAWT3daQHPLXImyR62+BngCZ5+F6oCnCQ32AyIOytrEGDt+DJh09k+Hd
KnxdsEXccIvFxUgPPllm3KC+HBa/+g72+X3lpiciqDzhkwZDwm/146LygMv5WCBAA54LpUqXZ9pb
rvdS92z2ft0Q8K5lvKfMfvSBQ9CT3Nn/ZYw6e/H8HI66FAfe8tJw+KesU1nHNu0QZg/+arlfYv0k
8j2yROTQLJ8ILoZcAysVi2M79PGWcMBvfAS3QLH3A66h1qWc6EDVOXnCpk7c3t+ctPDCy87/wDpP
coFtCagjoSHHR6BVaelbtivw3SaG66Fqso7MjBDADisPlmvr8hVhMmJMYWhO0zPTevZeXy6YaZRM
tf4n1do/hnAwUqSqAM1Bjrsk6ahHmbw3zFqFjkZOOD7GZar8rL4Twk1XeFs2fvDvvZp8mBTDYWwO
zbtmjuFvC61sZhiXuApPQfPQ5bMpbO5CavDLldxgd36qLVqfdoVveTBiqUdKNcNyPNPq2WGKrP+w
ajqZsUsXmEOwE5VPdu934PKswWj3CICms6P63NxNbu22MsXnfMAmpKGAwlqLjedS8BVgaDWQThjK
dDg7SAtuNxe4T6+nWtG0yenEY0rN8B8QC0ZPTtMprPWrVnF1H4gTwe9YWyl0XiPM7lQqazvdsxEg
GsCOwT2ueTNnJSeX20MnNv4EryHmLl8SMnJQwVgnBLZ1gFIuP6rXTCJMpMX2bZLDGPJe8L+QehvM
aGhjPSNUiOBh9v4u6Lsf6+xvsR+H3m+s36nnFUVV1dXREbR5nXtJ7NYxqf96LqvTwazLefRu1Wyz
sQcMTqG3BnwYkq1dOid9KnnJjc9FbwY5e4r0Bb5BoXPXokWzStm+voGSKt1wozJwYYflihbIxWn1
/mYqnuSVugjwgqgljJyOa8oyTz0Nq0CdGCOopzABO3Z+f6HvnEbnIRL4OX3h5FwDJeoP3tc3btZd
hEB6y1fueiG2WJ3V6WO8PNoZvxui6AEHgsNJBw+FPkTaiZT4oC4O7CgXTou+tVB15MofEb52vKZX
bwAd0oWDzN7uwYYwy0RSs7vS9+mIqwBynkcfGAZjENZIQ51Dl8QpGBtymXJ+Qe4vdQ3XBS/y+TL6
JevcWd1qJsMtF43IbpbJZjSSWEun2YIT6NO8obU067bbMvAdRIeBilDCdBO8S8HzDsHY/vISgJCc
gKeyo5qw5dzW+GPoCB0AB5ViRtjwndq/wiprlV0blqhXnq+6Xr4oNU8obOXxZKAUk97oF0HEqwDl
PhJrAaSCt1cujLVg+JGEIiirJsIFX/cKCV3XBIAnoRZ7BWg8uS4cSgcxJcH0FpHNRa0IcSYj4ccx
LRAWWfYCn4KzmBpJvop3NK6HyPi6XkCLHWm3C9ZtONN0iiCduapk63zCvLV/+FVaLtIAO4bnq8wI
hPqxm9q5r57YhzP870QGwPhUhFtgXK3DHRMpX0+/2LI0CmrPrd+Y4J3mBBAP6nMK/jp2WY8oYiHJ
lQ/9NQBp2+GhTuI0NytCgHdnM1w9w+fzrr/St2cDGriCcbKY3XCoSsi+uRibfgcRbl5j/VO2pIv4
ceykiU21Hu+O6/ds822jwZnj55Cxs7+upfUGb3CT2PylTg+Ne3XW7RjrGC2BzAtv+j9hoJznzmqO
F6DEpknSoLgpvzMYwOxa3Wp9AqQ/2qX+B5ZJQman0P6uyv1OLYcJEdvu/TAM6mfNT0GWtwLRroMU
EOHiJJ2CbfnRKqrI04n3AW6UybmvXEbwO/JYYxw+d5dRdldFcwnTaGq9SC16Ywm9pwwV48KP9t98
fazCEd77iRZV4ybbr1jr7/KOgUo1Yn2f5dQSdp1I1Qh+9ivA0fDQr4UjymAjoljmNOXcxpL7eH+J
cK6EtlQIHQoqxqcFnNraQLOstCuED/Nx33wGUcBBVRGAfdOy7fjRtGrihaIbl/lDKSFZGmCYlpEi
2TMskvl5j7TNI+DlUEXvuds8gdvkHBbIL4g1515ofnKeecQHO2pCpUaHdHaYFeXQpecuqJ1xHR7M
oMW5fgFJ+Li42DZXuj6aoN9H3HrZXNre97V9kmtep0rjH6H0yZz4byccg1apLG3F8BPELbIhxuXJ
JhcZCLTJPUuvXB3gJ8N2HBrAwoqW8vwjXXEaY86/ku50/oWzdcpfl3mAl1crjZWYJ6gU3lCaR+d+
TIQZgYrtmShMme1dXVH+fDUSwFAxQrGryGtk4y/Meg1jYyoAzvKrkz4KXMBlB2984x0JBGjVwfdZ
cCsqXaGmpxzbi5OYM3LsB89l1LzTP9OgGtgJ125AiDFhNQqtr8uQ+hiSLsUILz9uiRAidCm4+h2M
C1yK/GLPUzaT91jzbfO1a0nf/Z7H5Q2It57Pw4ay/+z+ftNrJpVSeR2kyVNTSAmKyTbKLBN5G9DU
FNlwbO/DX9yaG3bvxPFarpuMuR/9wWy2TDAB3H+g9WJUDCxPEyPTXGlfLgIUGOKkucLfaNozG0En
bRPM+05YcSElJqwvHZ+sxJNvK1ulZZwj8t2R/O2gZeC2ZHdQ67r5hnUlYz6JpXFEyC2UXsahq2Zm
IGVlSBP6ujHcvdV45cXviGEf794XPZdehNxQz5iX6hzvCuPEq3xczzfX61ZjeqUe0QHWLYoiv38r
6dxq5f3Rr9C1Ap0rpPAtJmkI+dbC3r6AaTHiDKgXoIDxAZqpM1A5AmPCZoB9sv9EAa1atNfVRCFN
ywi4fhnsD9gciycrUh30vVSLO4n0NdqOPNGjqM9+BluDTxzG/LrgnIS7URokMLw1QrtuEhdBf1bW
DQ3rMt9up0VDyD+4KQI16Xla3nBj6xeQWXDwKycE3rN45qny0rt4vTSisrZxcSsb5HGS197WCQy3
wSQub02G9awKp8Jtqycdy3EbzLpN0BSzyNHyQzHDYUy87/mX2clMg2sv3J5DzEBYaN7eAzq8cBsn
AGJwq5jY+ItREDPjJn0E0ZWHa8CXzzEqoVnv9J4LtGibOB9CdvlTY8M8zzyUdcHW5vwr1R1LcxrE
A1bnCW7rwZYFw0P9FlzElZfbvyx3NAnfi6mv4WFdCf0JrQrULogeVQ5N/q9+F4IMdCRXkRfHA46j
spW+ecE0X01z65QJmdi+Cqz3md4J+YOkqyK2ay9v+J3BmeqAlVlnnUgaE9VRItPSQ7wzOQUqyuQN
E0vhCRNmdts6iddLZZER84K8PZWHrpC0jCU608EyMS5eJR/5gBJowHu3kJs8f4PWbEqE40C5IRcz
Tr8LBI/OeIppZ6LsC21qKSkGfN0lOqifpIK38AEsM4xNmCHW7pQ5KnMMWKqzRzxHwAQRdzdZ5sNz
U85Zp0NW/mTki7PXglwGZ886VAFLeolBlEzemv1Gf+kAcMsAf94A+SrgcVQEwkInSaBm8oDT2LNj
PH9aBEQo/ftelpC/ly0Lp1N3i4wLyiXtvWWeJTiRYU9KO7O3/b6pMJfL5JmT1+NZ0CFeHI+bZtJO
WGpcH+R77wSU2lREivAafka+dgi99uSGgP02KRTIBdFm3dqYX+ysTXYfQt92k3guPDDyTNgNusGG
gLArCRRIzNxFsoqeM4yL09U4x+FqfXKMm+0CXZzNMKhxOKZnGNtJD5B0g2pRzwJzN2CdnMlT2yQZ
OW2/e3R3Gj/f0sdZmU9lZay72K8FE3bB3ci7f6T3jisnabmo/BfxViuz2r8asyQXuLZFY6W3pog6
AtfH9UpZjCahXAFiH/5DwvRnm+iauHkCBwaXovblFy0anO00T2d0mZhCrEo+v0EHFLh6ypyhJRzm
67Bj+CJgL11hPBYh/Un0qOzcUfCAfF/jB1dk0QrZfvkd5GG2W865KLe2jDhwANWJD8SMUtoV9BHa
RUeYE+1GP0TkPOM31pu7TsJzdvP+jhqrdIYPZELadRCJ8HcX2LG916QQ4o0ElqyOaPkqjB19Ji37
ZDq5lmWCVwgPRmwla7ehHzCZjYpv16veTrR1mZXgdnVU24zUQ9xCJHobPdmABHy+T7Z+U5oQayb8
PDe+jZR4gCW2ShYdbW5yZR6h+WN3fl5+VMmrNc3WAu3q0RaqoibhV7rPUyL+BPP2lRR53zqN5h8F
EP+qpAs2fD+7wAfZc97FXPl4u55lu4OQVcs+XBiLAx7f0aj3Ycr1dQhhGtJWqbaEHvvls9q/0e2T
rATizES+m9v4q34EAej9IAnznlFaly/yF48BdWa6+UuB0xuooV2K/YYvzvphCad1O+vNAonGWs8m
OOtbSy0iCls/f0LaHlc0Gnji8KH0fNrwIkjGn0HOc1NwjLWFc+SFckVQkhZB76qGNAheSQpAoKvv
lam1mJcNpqKrSHmuPRblPcixsRRhjKuHd3TTIrHmD2catJOrC5skha2OJ8YIYHWQPNxKTuYuiByz
B7Iuzji3241dxLzMVBcPG7iIB4fZMMBAnUcXXhSL0/bTWoz+W/Bf+gfLET58wloAulpQvvct+Re5
eqqEl9u7x2QXZzmG5K9zhfgWuCpkAHJXRvhcTTzu2Ujxj24iuskepy/BpgA3HjpIgB2xU9QcbXJV
eUH56rYa+sgQCfwkXeal56s60qycWd/OLz77ADr1BqyLjicDZrZWcR2ni0rybQr1+2p6/PcCNLTp
C74rsfIbmatZKK9Xxq7ROmh1cOp2Yzftu5Ujg/Kx68Ejyy46ai/7z/Vx1GGI4QAIiqjT9DZAGeba
ZjMysyN7cemT7wX7iKAutL1ljDVV2Ykoq/h00QJs7fCYIM9vhkx52Ue1MWDJlMMKr6m8sJ4hTl6g
4XIVhAMfghGoF/BeOzmnpXJ/1kZBJcx639IeSz29O6cBxGTqsmk50rF/WhU17TXUtHllg4HwFsdZ
TKOTWTSEPdMFoBC/rkuFHS4teSZ8qVJYqAN4RgITWAtppCtV+J2/fIvDjpmjyyqJdv7EALJTW+Kq
dulPZcqdRJjrEqgs8wRKJNNorytly8zypNrrzsMzZZfSOYgmtySVJp/cirZ/JvcQfl+tFHzA1fxC
6QgSlWRfY/L/RDfUK+yPnRvfVxpMEQ85s+yXU+rRwWTtqz8ntlE60Qv8ezcOt/A+mgDeXvqsJdVL
bkW8h5coTrdXjzpWWsX+XeV/tOReQw65uj+tUEC+Mjf2uftQbFyiT6ZBhW0+X68j9TJpjWCiv8BN
8xjJzIPbEPzpQZKNeHMMzhxyao4DqWUO3Y8GVsgOlnpOhZ7P2cg/HjgSicCK/9RjdxaPoib9/LrT
FuDC/q4WMTrv/2l6Xu7tMT+xIbr+qMv1brcpqdB8U1uElZYuPxEhnuwSxKbLqlKAHbUVl0kgODB1
MpQ9tjdalRilgybMS6Hg/g4OFruJxmoe78sEgSXgcnZZqxiUvACMeE8pFjuKlpekEuc4B2388udc
IyvrN1IQWy0BhuWzJXF5iLBvRER7FlnJMVD/KsSrY2goPSkb+zfsTZj3bkQi2BkTLWNA2TmWwkey
i9gfVIYn7BmGnyGbPAr/IKQau+4v3//cGkiBa9dwQ3pHsL6r0UJtatOPCJlQHbvUwhpId2oKfFaw
1Co/WK/skGel0xGk30fv4c0xg0kwfpJ5RJIb6xEKgyf7IMQvigGvU13qnzLrAO7pOemCP3tuPqtS
mp8M9uJeYu6XZLJLPNMdGEbKkwKaz9RgTfHAE9oNTe/+dntu+JGtJINvywy9k5zPesvpx0OEqMJZ
be4pRs5Iz5k0iZKmL2A2Mki0WZpO01yqkhHiRtQ4dOuR9tJk0fM3mZJwbYlFrXAweky+G2tOENtw
3VljLqN1KXma26UV/bxGiCYV8BnEPdR9nglblPpkBqDZj917kW5SG6KcrPkEFnWmNkBCvPHrq3DJ
M+d3go0Yoic64OKaxof53GpRQ89D4eIh28Q10k286WEMq3HuknysrLsij3TWNfMkTI1PSQKHkcN/
LWDKuGqxMiDvdsbwJxaePQ/2VeE0/wQzRebdWTtIDhM74P1io8EC4RQ2m7O+D18fDljT7pjA6Npt
yoGIMCiVYRzB4EGvTDzCvF3O7gkCz5zHRmBVFzafqV5xBPL+LCA7azWBIieecJBCj391aWVNFXV2
E7exan3Dew69+MnAOR5lek+WKPgwRMogOYdrAbysKNH40VCLzLPM9ZTw6migGxSFXjht45rxHwMQ
HDXsV/ZRVVtgDwTxQXi9joWsECeZ5vMtj7X5YM0fnqUwKbgXp/+3hVq1f8kkS1tDdzwQrHfOg8tc
7jKFvkH59QuyITqcTzstbTFU4DDAtMqKEcVc39tIRNu9CQnyww3uU/8JKBNx45o3MteM+Ct5F3Oi
lePnqjRzr107E4ursXsT1BrTJL7gJVRLuEMyGGhsRw/m/0P12an7uIRt7gzFHcrjo/DbFVIfXhS9
36jB78u1qmPhz0mnZyYBOBivCeukYOHripkbIwTPhAxyYl7ZQO6aPwPLip1RX8ChFadbYl44Jt+a
Acwb0LbzneqyUS+BJQMGN13OX1YWvS4xqTjG3jbJOGp/+no169bL3HCJysWBwC6WQhgob6rr1gj3
ZEc1j1+LWDNO1Q31qiBXumEvYr27TbCzo+VP1X6BHIbAWNS7bhfGO7l2WoJlJ7eecsSvyTepavqq
XzupFCf/IzUKjyoXD3f4Ttdy2bdP/raaor6iocTbyYi5lS+rrT5K2ZS8ZGBEEQkgMdHOBUbJ33Hy
facV/ajVdwB25S4PQ2/r3m3C2ARkPXbmCm2+OlbkJwApnMM2tM2giENb4DSE6g/V4OxL8xMSo5my
SDLajeyaYUHT1T1DLVO7kq+UPicAj8/Gy54GvMRDhcCwbqyvFubjlcXj6rGkx/PzICqddy4Yt6ql
ad+2tWFIHX6WrUm7Nvm8vKDu02ztCsS8waD2/931bzoQWIIE4LtGnUz1UjqqYK9kP7eEmbFEdLbQ
vC2VxqHfKJs9p2wR+V+Z/ueLGkWUpzqXcAvPTAEEHn7eNPVmPAhBjw2GI3y9BBQH9c2Y1/U86MRT
VmMMFyRexWyJrZ+1R8XEsDRoG9rXINe5/gsWDFFpH9TwxBXwDeZzf/Mlyj4E1zArAFrJDrQuGIbf
eQYoMm0QW4ZXB3yIZODNz/tYziU7QC/o+LjM89W7/7/O75x+95HeH0FEd34cNBLiapIA0kjRCY4u
XVCMFuxTCN5H7B3hjMvxsjoiarfKN2qGr/k0ps+PO02yh7BsOswpTI/vr3H4qnNfv9hPC4RZGB0l
ERSDqkCdAevPoau9jTfHFPiTkPcGNw6y+V9W5zVVks2kDMeXUxZj+sYBXknc8U5Ulh6EqBatO/OS
ist6z3V6eXOW1K5H4+Fl5K/bgo7/0hTcvGrBTPJaE15RBk4HISJ3iD99Y66S1GFOAkzGv+3Z+9sb
LAIOQF4XE5nAZybvQvImKmbyIR/mbQXmpCnwVPfQkHsR/7kuRGDIGHWmGXO7VLoZeGJohJVCHRHn
SOzskn1yBLExkLc7VCaP3nwgdKavHEI4g5vnP6pdQS7sW0atz7kBklza/bzX/Xry1+3NC/yBIfDs
31l/W6Iygd7L9hzwWFAybArgPvFli3Sn5jNXCtuwkq62EA5uetUJM1ZgYWc6E4IpL3Uc1jUaAtTO
NfBOWpPLh2gh2Y1DmhJw/p3/j0KcbV8FrMAH93sKRs9PNFbPVwsF7XOb3wmcDohsckfBUKXMf8X6
UCjiYuY6oVYWaHuCWwqLA6e1Y2RMor35C1i/esM5eXvwr6d4AzGSRj2TZa9jAlt99tXUJf05I9f2
5Dw4W7rYib1Z1/GehdlMCTyHkybT15KA7P/WFG0ncbtZmXyPj7op89xpBIdz2xTHiffIOIQbybaC
ZGL4iUzuHbF1UUS11HoXPdnfqVo8sGtQxO5fHc5KM43fBLeXNhXuWH5IT5oBWXLisg1aSjktPv9j
a2tTfsyGxxQccyV/Hjiv1+FKW3/mvDx36FiJosej3b2ltX8DAJRfcNyf9hAr5VY11HLbKhyG8jwn
wgDQlAT7US8xp+s9OiWHo8jdADt/Ze172yOH4WUWtc1qKaL0vRfylcA5kW6Bf+2X1bNw3xDNxRsD
JwxVmckUfIbiMAqVZBQ9R8GDXCgF+3Xm0VBDWMCo0sVlibIly6a/PjELFwJq7xWz+KH9h6yJVYCo
NvEqYQUXHItn5eq9cRXvcdGnhkq5YZ6Hw0I/h2f6ebacvPcfnBercYN9RVxhGA9smyquhVPbUh/X
ZIm8pwMtomHHWyo9fAY/QJESxD1zPLn1X30n1bqam3zOqGsI9HfuEDCkvWJu9c/G3fzHuOqOCiwC
z4P4U38+rCvEwrCuhiRxsHJyv8hZKsz069/1o0jEMtUwcNBMQZNG7dpZQkfRcQwpNW+W2/np8y2m
7QB0eM8wa+CvtyIq4JGHP7pEcZ/PExcYCWO7zjgi8/pTvVQYNu5qwacgOWgpVIFcgCyyst5tl5OW
kClZny2qNdTSAL/IswMxR2evhDjeKrohuoEw7kOlIA8P23aAb/hRNtDHVLGUdw2m5Szc8O5a1QRD
6IZ7oqJIwI24mOoMhhDDTy3A4r4emKqvLPqqskYnjKjsYY3TFkJANktrjuUcxs7aOBZLQ+7Tliff
6pnrUBwz8N+eS8X6oxFlv2ExIYRE58jCoYalb8lw/C2cp+8WBo0a38TovdyNZUiGlcIHv6kmjpLx
eI8yXNjV5MgKCr0YhB2os7nLV7/m9RpxmRMse6xqNCRLrIeclGc7ugCF9v+QenAJYeG72+j23mRm
E2XTQhVGW5OQ8QLX3rnozhzIctAKKLKpV51rUmPCVNdRMw9s6JqgT06AcxLtOdpS9BCxMqIWH4D+
MZCvMBOlKWuSU5Nv/bJRKvpVxQo6VJzEiQbgeabFHBAHhV8xLT4ckOZx6lg5A4/l8ksX+8TL47Je
GDjSAoM1x/Ytrv95wEe4O3FCEc2CrXd0gmjN9Us4fW7lqouMl+B9ScAama5Kw2F9MdeEdeULIYvH
AiZuNQQ0jr4Tb0yJcDE5FWtmggKiUUvP8NAQO6I8BmRzU8rmTslfDJ3kRjDmSElFxLYOshUUuI58
5vzUDhUfjXNv1c8h9WkiX+4BbZD4XxCO5YwikrW/Ac0TjSKSLLqkQ7ZDNKAyXJoStZR9wSQ709KY
/AkokDv3HlU7la0fKfKecrX0xvm+KZ2Ng0ID52f2c80QPECGqUn7T3H+JUqG8zaT2LBRdJl90aNk
QDEP8Iv7iY7BsN6KFFfj0fNT/RtB4UspP3GC6fnhQk4m6J0oMqgdTbbepMolQ2e5jmialCmP92rd
aY1m89bj3MjbnaXxQ151DrWH6KCsaQ1Jb2X6eR2Iw25/tVcCKOYeWEBLGs4wVBGJcOGgtcLNvH9y
c2mFA3zVjXAEGHS+J2vKPsjVIIkt4FtfXjDrm05VUbLTr04Hj8pnfYmktDMTrRQPL9GMM+AuXJJM
5kvaMPgGZt7AyxjenwjVxM5Y7BMubor6HniX8hqw2jrhfHi98eZEbBGQ4IqjcX2RS9youi64dlI5
+ffG618jo99HKDhQM0v5LFT16JTx05Uv8F+quHKHWH9D4ny4mzoclFeHQW6GdaMhPUWMN05APXXc
Q32U3VM553yZOHlQs85MihPDYT8ayUmwwm+jW9ppGfltLUhM7ku04KjIZwWPELQ7wRpX3lkjWf0Z
l8usCbBaX90/SsKEp2Iigz19l3kJJIBkU98ThHhd01ypkkzgEUovDfULWCL8e8dSsW4HTR0rmobJ
OBmlZrl6LgSIS1EmBw9E6yC3zcaq/kAaAFJVpaAEyITmR3cZwUHrkCGnLBQvDmd9d3sfIcHNVHkv
7m9qPw8nYzydgxdRhW94mbSLkxAJCVNq4YZdopNRr7hWM7Tovgpr4d3zdTUbSd8wHZAeFA2p63mM
MKb52nGT5jZDUI8MbY3dgGyK8DLW0rtXUifOf0rjPg0gWpI0tcvT5up0zP+BLz/hKYc/TbCBsN0b
4dy66Py1RGW3bXIgqxwuV6QY42sz8M+mpw2ry7J8mK6Aest8eWqsd0TpSmrgK7eE4QQDHS/p/wt1
Hq7rdE88s48O248jSZxPC/Oe43IkWg1N+07+qfBQnxHJW/YVek4s7CxuaEEy2RFHXdytyihBA/8l
kGnUzKErRhVwrRPh+gVoUPsP95XV+ZoCL8z0IXySnK+Xc4MwBsg5aFy/eiCdF7K0nulle/TQoOg1
81aS+fx+jDqLGDDF0a7kE+c4grEL4z5Ao+LEbYJ5KP521XFgzHjrP/6anwO7RvEgIPazFVfn9Q1H
n7llhOtsHhioZowecYoHOWIswxHFSkElC24PJDgYrtEFfRBPcts2dJaEnlAFwThXqnuMTQSRfisM
4QwagtaadOPEcwhFrgHe3aa7UDp1D84LSYTe/WEljAm8L4LnGlc2sxVKzDKXC2Yi6vOjjDjuO4JV
EwNN3dkOAsS5Fei2XZjh311j+qqsaH8CbmwrLMRzcxWOvX1xLJmtdkoHp7CWeW/i9cz28Wvg5CRJ
s0e5+0fqghru8+3mkIZ2OEe7/44YHDO0mk5r0o65YMBHlzQql/Em4NOigGuGt0CalUUQds6pLobk
DWSasuQK21xa4YZMZZar0rFAmEw40mN6tV2vujWk8rZAOBzO3ywPf1RuIMoDDNURKK46RJYLAk1u
jYMeaXKDWHmx74hpeIJAB0jspWC/E7wdwdMmEOr+TFCUnVKVvjA3lTHgBoxqOgXcjFbPBb260Yup
BjB7I26qF7FjuNrv98jlCpeS9h0VahqW0bXkn74sUtUzAPo5b1n8em72w+2Gq0++asQJThFqkPUk
oS06Fe2+LzI2moOEElZKXPC99nzhLpBfuNrGZ6KyoKsVVT9GkTUB/qvYO143yGL8QymHSCaowt10
3R9yDqIgq+4fmOa7YUIhpin9rt+cMM1th8XfuHmkdcmLXpEaZGJppig0MKqX3K64HLcNtHAin14Q
Nj0kbcQHouOoXoIEYxwJ2yqre1lHj5NOrjkFe65dMrqs5+TC/szLKwTY7BqztERZJecCQopUtO2e
SMK8TXjLwVRIFMaugKXTLKvcO4MOx0BM1vvXAQVyymTPJZ/ompdjhSGOiaMPQiosfTKJtRgq7boh
V6GML+fXt2ncYBG2ys1uvKuEtW2XXBIw4+LhEE1GGf72gkR5qBoa7zykuv2EYdjE+vPhTDvmJN77
GQUVKQIm0xYJZHWjDRo4DyV+ekNyaK6uHebZQaNfYHTC/Dv7rEONvKyaFsbFsqn7F7tw4ri6pSBY
gbuTuI2F5dj4gmyupcqiGt8tnXgu7eAN1b/cTjN9F09hU/AXHV8IlAdzGnfilPIXgX1BhgjWMpHJ
wOP8XNuuELlZLwpX8LxkiSu5qZ88ReUfRVgvhSHifTp2AHwC0DbWLKBoeudk4ycQJ+nCv8T+pqEa
p9vuOrtS9VdW5xS+wtud39AfN0wzC+6qFkKqEoVoeLf60DDo0c6ajl5HU4DnUbcY3vxpNgMkUPT4
AFOIyvmVTbS4StrQp+xZumz4k253CTHTtJX7qYbe/2RxvOHXsqAouduVTNvJyv1/5twPM8nEwGgz
5G3NGTexXfOPVBN85A31xAY+zdP6VC91yhaxu9PJbmizJWMwZ1/3DcLiXAhTqeId9p1tYuH8oZ8R
9TOpLX5h9JTkZU/17ox0XX9oD7tuPrUR3xuAvoTRxuIb1x8px+TyJ1KcTTnVAqbFNx3DE82zxApQ
d2oovKrpFlVgHo9W0dSPnb/UZCdIBB2PREIlQfy9WbUegkNCyAjCdrsO0AnWQcjGN4GyytGbQY2p
GOknftdUaLZg56YLr1l4Pxvpr4N5jDcwwHZgm6sofvvULXpromMk4pGuZ2IXuwwxGpjsGIimLQ/y
Wuhd9M748FYwzXVV6JCce66gAndsWCq6a5MC8a5YtA5ONNkfpynIEtBZkyMeSVTgS5v7oIyEvw1t
ph/gqLp2Z8pbYbPeBHWBOlgzzU2PhZwdQWZBPzrIIVjU6O6uyXuwzvyG7OPIcn7NPXgJUsqKJbjr
ijZbvtE/FSUJivynbHpj99UG4JHcsRUiwVIWO9ySjat6t5YBg7WmQX8FfcJFPLHo+ExNgm6bWQOe
ngeAJrv+NDXyg97e6GQhZ6cYltWTNyZxvME17Epy9Ar7pKhCTtEiQST+VGSohW0jUtg45mV+oI9X
X6FzRGqLkNg9bLzoujQwDAAoOAVwYHGBJv4m6E/OfSc5vZpE/Yk84yTY0DBVNV3yIBaaCyXKyKB6
wtsfcb7QShv/Tm1ED9lQ1KMYMXUgRlFdQv+sX6LTJwC1VnA8qKUr67by97LmcI7kjGONscOJGrwX
+rl5nfopKol2K3JI35kCP5G1Xq0t8ki9DH+SIUX3V6/sTsyPqiucwhhVGQK6VFRQtBmQ6uGgeesn
xFItTn41Ala+AzEe46CjzkLm+K5gOC8/a0/pdKfg1zD8uoLQPBcxIhGYC2O/sHBc7AdV128BioBT
l9iJNGN1hIuIEG4kQKlNvMjyFFvsflodjNKaHAWF0x9BY43w45XM7OxjSwDpTIDZvt/sQZF0v4Pl
J4YvuJdScZhFXZ+5b5hZWUxAvCFnt7c6/WFaAgWZL72xoKXQIyI/8PhWr4U2rZEc1u9jPoyicukY
5RucWjTc+CCGzJE72i9tNuIIWP70eDmzCB8Uh2+r/DeS78zL9abn60F9QvVvHklSFBU6z5fi8bL2
W6B5JS9EEZHKXFxhOkl0xHyoY6krg/ita1ANI6QAc/s9jqsCv9sF+rqcqADMZAeEH4GmTfmdgZRS
+kH691r1rysCuXxdGNq8WoE20BHyUfGlVoXkDeIL/qFcgEWOnvGzi35pmzTWNvvVdH5+J0fzZmr3
bjBe74Y+QayI6EEj5Exf+H3zfo21YPcrPlIul0T+n+2pQywWLsBZGTjErcrKxbt3eGKsRG/GzrKe
RLcQbwshSH181DKRhuObJUjaMPLFHHPeFMe7RQDGLVKf6DApJWdhZ3MKZu6jGAW8CTGH+HUTsZu0
XVSPH8bPux4J7TN8qvqQC1uleC6e1/FVfvaYYjFaPB9QMNIujrzFbtd1LAn3TAGsa3qi0RBYetwS
/S31mDBYjsA+1KZLmR2fQWeK3Y91VFyGomAecYM1EWkgpaXVWjHrLpZyO0Wr0oEflo+AuJjF10ws
EGcaayPIT9NmM83LnQIgNXFG5wmZK74m45vwC+S2kezCT+HMfRGi7sSeJx4j8E8m2ttf/3muTv+9
nDF5rEQb7mGmIq90adeBpEUZ3GvKbxqFQkD3rtTClsvUt24zCyZG4yTUn+9p6BWhJnF6udgwlZ5D
P8g7boIfEmh73LE+IVDIpgiMkpyHm3i7vYUtge/Tvj0R6vxK2+s7mLZuM5d4yrlFVksuF5YhUyfZ
HVP2QnsXyODkLGGDIfUEw20YXpmeZy20Il1Z783FuebY5WeZbCcQKWXg1w99qNgLf6nnostr3KqW
ejwWhyKNOG/+ZkspMbl6ohhwxu9PJHKgIhNbpR3a1HHceVsaHFI7X1SKEK8J792Od99dN9pLmMlZ
h+JD/rQTJB10+felrX9mu2arCmAbuUpb8VJVK6TS5g5KWYvzpHE9FsyFDpb2ryKtRhl9+S78bSN4
Pco6JCLj0YvliKkdZX0sCYQrsdIh8PFUz0xrTBJ4sxydnDyVuUQ2Lt7pl/C7Cku1Vmdz1zJ1ZM/v
aBYTARs7C+yZTi8vmimMHM5Cs0hF4hFV1KWApbWXxLapDxhxdcfl/xV9FZ6NNEXMIBg+BAuvLPQ2
ZDhHgt815HOP3ga4xn4JaBQsmyh7t0FVus3TzUpjohYeRrbKTgugNNxscuCakVh9ar7ZO0httDSs
5SExzJ9PllAc+6jvQltxhWCJI3nSuZx+HzIe1AymX2USITkgyeUFBUpvRbeS+ZrJrozz8sqU35DG
cvZYmpI6tujWNl9ClcXIf46vL9EPWINbvwVqSgl/fYpQLl0uE/7zN85Y83veR9Tyu83T//GCW9b2
/VlL/GtGgBX8z3zwjxQunbVdwuS5dt37D6vb0qCx2SdNdl2IYdqtDi8Jr4tTiKXqJitb8hLwkHpU
+5RjWmO4TCYWJOPV28xMe0/uffNxzX3HUsLD/WVntyNuuk6N53C+CAG+7AGihjiFjQYuVGBjjJ5L
JUXvzHSH3PziqLbn+DF8A9AUEFVBidJpdvk5AEXBMUbIi4OZP/m2IBr4PbsssEWVxG4SxPwWu9cs
8v+uU1L8uduo48jduJ4dnsyon242cRa/lnPs5hOopOiFn2+DWxSvHYP8aLYtO/tbxeOlvaFsm68H
IU5Kr9eKdeg9FEXvKT8DjUxh6pW+PyRh8xKkzrcyiSL6osZUTL/mfoa33CqW/x4lMwgQXlcrPAX+
/EJaI82aosfuvmt3SOT59A17m2dpmJm8DOmIdDKm8fpPh8Z18DN/bcGutt10ok4+N2weev1ZOgG2
91ZS9aMZCEWwjUII5TKTjaXgBQSiVqtJAP5N1MUXOoTA7vp/iSlMbm89kbNqsxhH4bZlOxf9x8wY
yiE0KnaX5AbzGX6ZwSrD7cbRwe3HGrg9nnrQ6VBcTJA9jpUS/YYV+8gVhfgfJ0m5X4SrIRVEfweW
TcEIxIMSvqhR3/XIQVNdqsGuADeP72sok9UYIV6flu07Kci1P3rZRTunLP0+DS4ouLKLuKcPZwOC
zuVhPpBrNyhLOxwcBUc2IEMvzkZTYPz1tMqKjxi+ZKxqSe38m6Lqa5fBTnIE8T6V11ybrNFHm5wp
fRY+xxS2GhkckdO+bgT3yvKH5wAeV3wb4q+Xkfv5xFAJxmQr0qz2L4BH1sJbm6fpeXw4W6JqqrlL
RGjUEqdCJWbvqzUAGBI5ismY/EfxvemJcbPlcYDZPenxdpPT1AyV+qo8yrBE5HIkth9iARWU1vVB
esrJuHMdtXn2T/odou3opN1UmvtLOXMSUc4KFi0gkyi1kKFnb/i0N+lLKPxzC0W1oa6XIkb5xnil
oTEo2vLp4jjLeLdUXNkEOF1QSK3FheWrol5F+Hv7OXrnIZnVdOiPYvI32B3rAO1iOhEnqGc+epvR
sMHBVJ5hdVySman7vF1RXJAm1DLkBCw1s1pmKPv6SkiFWDii0OjwWd4rPBLyrtAaBTAtEIn6mmhp
X/CeUQiKM2K8d3m+mxljoLXQEkqpLOpIIi6hhcEejlznzeT3w5Em+8LEsyPrL7KDJObdfIhbrS0B
d1QkE+5widHecw+cBAsoVXCv0Ut2jCOlegGBqCktCVj6yak2VRQeWW1CW2NmaUrN3ZbKJoHx0f99
bM28S46UrikKZjm6USixNHL7dgk9uE+fRD/K5C8TA9sEwBFB+Jom2cDu4olzRzlHNQ9I1iZ1cBfu
CCC+8+rQq8KhXnwPDGzmMiuSgGVbeNmC1Zirq8MSyXosUXELqbaOpzeH97hymw4WiNMFn9o3UuiI
gbrRSnxcQN1BSTxl9lUKLfn3JG/wbgmAJZqe0/KpnZTtRr1fmJZ3Z5kM8KCS53D+6rbZgWrAijTd
aVRIWDTibPVm12t+1t5utERG0tqDhxQOJWPTRcfo2FCfDiXpzse2cKoTasrqXm91X6zWg5Ftu9YL
j/qcxvVCBCCchjUMxlNtWJU3rn30P7aH/geiaFaTEZPrwBbHQSDUU/aTzUfzVr3Qt0P1s20A6Kpb
ZEYjbzV6p5pQ/deIsiYGPLIuenGtPcauEV+nQi6kxtKFlT80yRAKuGL7r4YYzIMtndb/VPriiDle
PKxouj4W0+LYMmi/iwtgzPWEEixF7ShgJSjBP7IzKIIgFSpqk7dtTgCNzUtxv6wSYn+pulfn1E9c
TjgAxlrNwH4hbbZP1Ukb/Un8QxthCll0MebU7BIetCD9cUj7HvGA15lOzQhE8FRewR+KMQsF67C2
Gxz+2lJh/Sbckft86MFfl+hGqVbDCo4RcNiYF0a6V5D9v7obnACuy+djl4qvBDJOmDWgKLJAPWqY
7yxxEBnfY0Hk9fQVePzUfnTu5V8fDWgutw0X/S2piaLKflOrWIjvombUiTQZt4dQAe/kwnWkAfJC
Z8X3gagc3JVbDzK2m9eyWWyugvn6LAu/fAz/4l/WXMXI/0civ0lHa6Acx/ZNRkAQo6cEbWkDoFtY
cetW6/QWceWa5TRzfPuDSthEBTNtGpOu8MOHmzQbl+Jzl64k8XLxkEyD0zuznfSD3nCc740VAQ++
pebaoAX4t43keQ9nxK5b9XHpFz/qos5QIssrW9l2ukQlRz0YacHthHpSd+0COni0G0DDiBn5jb1p
0qKydymXWVPkpaPEn9ot+VrDCABV5XUEUSr+tCSKlbmCU8AVfU28W3KEGMT0emF10dGnWD/tTaCg
XfXDySBoW9iqeu2jiqGvzAdvHQq7HChZXqVNqrDdtq25FmvPyYjmsxpAHXmvvWmQ8Vm9zCvDnIuf
Qaz5y7h7HCEhH3M9bCUZw6zOGhwf1lDKwyAuDDLaXLzSVJAbfjppPSidkJUaUjLwEauDdI5GebD+
sAS6189ks0HmvcNBRghO+x8mJX0vNtsXUErfZaqYmfZb27iVdY3AA1T4T5RypccR3vdfttPQk3M4
f3svPyMQ7/AP6mEOyeghuWshRKTVM4QSSIS5h6ag2PCtnxmq7e8daW7/4tvihEVN7IhCFaJuAFrK
L0EB5zoqIpVm7AcZNSd3aFfsWk8iNHj3noSDdmKg8ehCNPUbvmy7XCGaNfEhfgfD0KEpqwKMar9T
pUcGJkQP94Ci8QWB5VhZ5o84KZDr70Rn5/OlJ5qeRAqXCYxAUTjZHCnYyssbqGKGhcUF965TW1Xv
f7yQ90ObekTWlH8DqND72WxISYdkzYBqZ8uDjKNEHqxMRwIeT+Snlb+aefX2RnmJnsM3NFySNYuy
9JhB5uJ7q3Od1HYhHP5+6t7YACBZ1DqzaEW1GLNxKb8CXRYDHaCwyPQTcO38Kug56ao4PtEy6VX+
2izXerNo6GLuHLsKXczkiGxxSquCtafeNX+RBXhEo0v9AGgXCHB+F/gyTolEZ5jkaXwh8Rr8Dt2L
gdDY3iD2oz6nIaku/Uo9Ky2aEAk9vGFFrUCrAk/LcLqx5sG6uwB0PXJlLA2FdKOTHg3wgaZu9uJz
hdh1SypRCVZPcvG33r0jNnYvXw5Y8e1Jg7iunOcdZ47YXf2bjqKYP24zBwbgS90HyqgtYsAntopO
9yATOWDCvBvv4gUhvjUeq0QaO+LnDtpawmPd5e0wunijNAMVr/Y6Cm96OvCps/QOI15tz1uTI5cX
+UjbNSTXLblr9N6Ftmq6kbs6EsWkT7ck8hfB0PL/LAw0Pospxsrk+dpLBfUziCu6xpDqQOyu7JQR
KOxWOQQOyyU77RBRi/5PYvURJ1zOMhhXmoCo9vMAW1S0c4MeRFkngMpwyzOELCj9kedwNLgq8/Gw
S0/t9S8Jv27epOS+CTxiri5P60muptcwNp41t/w0uBNsyNFhkuCH8l6nw2R0JnXzmDiPv5NDn+SP
N7nfGfCA7qK3UlnNzxmHCkZOsZbX7rTuqZlLWp6Ytkk7twLvPxHBzjZ7AETmsyvIudxCjUHZjAuB
WZK5Ek7VBRmwhom+6LVx0BFAkyzMSh/lJfJYdaGgHFVlfHNjzc4mM5x8tZIsvL+OCc7ngmANlHpE
9BJpwklJ+/OSRpcT6bq4PUC0UhhbhnBQ6CUv48YvRLmmjhrI2wau6WzJEDnIckdSQETyJk8Gc5JY
A2rb7IQaIRkMmPj8HrSm9GnHt1mfGbZX+O37oY1MpMtiVH37Q/f3vUo7QWQHV4ZTOwitPto3gVgN
DAakA2FOumUhqlp3RHQWmeOULjGbaugzKG4D8T2rgmGb1pAZsZ/wX466AQOJkGFCzS58l+474/yI
1fHFkKxpg/0mwbqnPt4SNHBgsAJKJtpuSa/fvN9+0tfjrTfIXlk95g9xh+j/6Mnl5yALF4hQaYRU
XgecmoHAVVY85wq9XTrqjKJWa/15DuGbuBNC0i0xoxV0hfUEyYAVNUJt4IqyOZgLCQKCrVNu1v31
HhrYWmuxdteFjtYOduUI11/RQ+Ui5SRxXrAbCl7hccR5nDxsK/0aYYdy6B4qaI1I44I3crJsOlzr
U4Ue5G5bX+uEESxpJ9d37k+caGnn4zJkwTb7UldxIe6vHc3YXVxPvHNtoh0oK4butkZZgv+qM7nL
F28v1BTIuenfFjgZTbGgWaMhP8xLyrItUAO7t1hqGu3p/UjBOAZwsKpX7lLGC8kYZlnlRmnsjP01
hyRrfxIQjuvzOvkOw9zdfxK58jrl3R1m6IuPvrhbeZ2iL2x6q2JZsIqpSilUflJiQRVXUVw0GAj6
jn3GVcBA5A0hDAjF6Pko5YKir/XNtWUxJrBxHdWjETB+Mec1EI0ZNSTeqfx0UyrJDP3xyKCG+jG2
dRMccIS8jG4yxemJuidftoNh7L4puwvH5OYYzDvpyAwZLkzVetvY2C6ZS/iZkNE2f324whI24maD
rfkNoWBmjAVxXFlkDfOeBe87VrCCvZtRF3VTaH0QLZu9LiqFfolNKYnbOrgr3n47RyFvXUpetoMd
iksIiwcYV/WkdJhuUMYij09zGONeso0kl/DrqIYemJBlXiwz5TQBbXnYpdiBuuaVFwFR2nBQy35C
8gyMJKnrIelgL8phYo3E3Eh5x2EZQpEk+JV/OcRdMbwRYawf7441QzHLHzpALKPRzQjCwPV5fa7E
k7c8Cqmu5fd3jxU2LMOWCLiP9a2mgfUjz3w6gMljt17pV7Nt+VJqKWQIapeqt1D3pQcS5DwLuiqV
IR0gZXHW8X5ChVtYhnmBCm0HKXtAhPkqnTz56NiCn5qOdzhO7/xgVtgPWnIJNaSSsAh29k8eJy6p
t4Ozok39WvDd5OhYj9gj1gFfr4fLa6HYDqMOd29bPGIHbH3j3JHucfVAabURSCqRXDQS2O3FDTtx
TdZSyUABO9tEsM9aSgtvllQSCmN3RB+NNxfpCH9eqBXEfjUACwV4K92JatR+o0+TK2M4uYQdH9BH
IpmhUb27r85U/kz7zA8RyfYDBji+ZI9eo9cENM58K5YJsM+T0OSAdMIvDoaX9Xf7VsiUbJUqSTEL
7wKZPUBOSpmtLvYJMd6CwsBC7rmekeAnH3vhKkdQdQU6PtToM8tdY8S3qo62+lfbmZCLox47kM07
ytaXyN81nSqKefT6WzV1LgoOaz+lMjlpI3ml0+8k/XGHCKuR1RRUM8BqCDcTmUUIWNM1l99mNs0W
5APsservoxo/hI/+gx8Tchx9Zo8s6O+NrgP6ETDRMQfwu1NuJtypWrJ3kieoRLOS1JKgRXn/wYTP
o7wctYF4QL7yRCLFlwEtep7JmWr9R364YLNRa6H+97r+k/wNedKRjSVGXg0D+T+mij3VuV1lvqeg
4bGe0UNOPr4Ks7dGt5/w3m5H0qxcizaZ+pqeSC4I8/XWy7pE+FoX3g/mP2D3kSx4aRRT7Egxuhk2
XzivhRsHp7klMzyPCJNxeiL3khzr7mdkMRAT9MEQroSio+6r1cbj5p2QrbhSSMYUmJNDijo59DUs
+d2puCnWmXl24qYYx3kqU50V7ANkCOfnRztfuIFuvPAsr/qNJTnJWrAiTKjRgOwqx/HjDL6aJACK
KJ0LoEI0OQtyl0AGny5prCJcqUv43pyhD/9KOqHUQWrlWZ/pBv6pPc7OuZa+3D97fOi1EG3kYOdy
RsR2hLdX9K1J/Ariiig2DSOQgu+JnAcvf/AXuYih0kp8zX3rM687Vunn6LtDu0fU5HntRaFed4yz
Zt9zo6P46IZeoG/QigeLOZQ3z9cn5iIB9m4Hx7ZEUtMLQl9sBJZLx6ndeBjsVZshi8vGfyix8qQd
Oh5k69sVjNl6VeKyLYtm0LxQcF+4NI4MrsdBogmoT4JG03vxHl9vGlKH+gx9ZjRMlTg6/atRrEbO
CmhT26ida+WRILQIFYTyNGTmcAAj1BiSa6KhJn6cHcE+Q20GhZS4yOseL3lt9d6dndrZQ8VeKFaF
XEkRFtW2MKp97vlWFYHj+sEXxPTCVOgcvO6izOp5xRzVxYbcVZ/WOBpLVLqhO2w+hWyYARE69gR2
XpkCuIavZlgt5lLp5QnAM9uU8AkexTQtKB/vZrGzee59rArw9ufIW2dIkzLiKRlrq/sQJ6EhmpOF
tPjeumVxAjckg0NmwgHlUFtP/J1Xgwejk/1fOoqqPeBrsWkIqo8czTWQRUvsJ9tGC6tM8+FqMje5
GeQtBl5E7+lVmTGkiC5M2o+2n/YWRTjU8b5Q7YTI9NNPfQfh/pW3KeoOYTOTYiMTf2C+344V2Lcv
HEu2klVklTTAbWlqwbqVbt8aChSQlXVNSqFQdto2wGNL78st1Ql+A3ne2OpW/n3KT8f5iUdqJT7J
MgJuTpeJQLibLJ806+E8NYpwFzrPw3fRfpg7ghW5FqnNPp4ewlo5/LvNgTKSU2US8EPOvJBnCRPO
cN2SwsmQnWtIxnYYE8bVdh4Ydt0TEi/LpGiqHhDvf0gbXm5OYPRRCgurWxiyjENxtM2vjr76be/Q
Fp4nBd0fEwaa0mn7ru/IOvxdZzLpNGdP0qP66YoV/bsxNE08FKaIQeF2dgxJfFbGNhfHHX9txA0Z
ceGgKGR3KhGUM1TIoPZh8RhKgjmwJxwHGmYP8JasNy9U69gP6QZCET6nJkLfaEGHZc0mig6sW6+W
m8nJbehh0kBnqRxfogW8eeB2I5vr0jfFVoW8GRj/bXBTlsjDH58pJniwKx4pUbAHCS05UBHK9D4X
w+qDjClSaByh8q4qL5s7KsxSXprlTEHk5uoYBecY55s3jUyjCdr61OhAVXU0TzXpvtjLP9A07ymq
OykDW6/M+2REKoRfkT5arVQ32QEoswOQ9qudL7zRl+3dsMHvLm+WNS5WqwdAIi3M03R/Kr4V6dBa
aT1upAl+kzYx/B3NdiacQ4wlWfxD+Ji3lzOJu7oRdL5E0vDsKzRe/Lv6wJrruLesGVHWPq72SHEz
vlzlQKsBm1mZFlQjc99lIlusErARgP7mNxtW85S32/2xol2HcPX56AojnzLpjoJX9+/QpaNn70/U
6wxNaFYgsrw/dX1xeVKyUFuwPHIyK+I/VXG1y8wv5DmEJ6qh8lh4R7MQRowFZAVx3zUUnW4L99ER
5CK5iqSlS+AE70KUTEZkRBjk9Y0sQ4YrTLO+aQwvQ1fvy4325g0/exwVcSdm9QIsCr2h5waL34Mj
N+Ce6bOPVXzJ2P2eYXT27e6w+MuEDZhbvTNmMeqMUdOY/przxG8yxVbqKXRyYfVJTm28WGWeuXB2
4kqUFSByqP046upn9moiPt9HJcQaRo5PSLgNru15XUFkAOJSFdr5jFpQK7UhHRDTFEHxxVkZtrAl
9HM/kx8FPnjsOM+ctu8s7usPeS8ELpv+yFIxWd2OA06Vhr+TAu+Gx8aeKF/qlkrzmQ8J1Rs5rmdR
qBmFd8o3Eo6HD1V+s+BK1AJpv2VhVRa1B9Ukzx5LnX8anNwIyAxB8dFSTykMGJI1khZ9yLd4oSDL
L7uSlmp0ZvYo/6Y1zyoJAluA+uNpA6ZZ2D83PYdaImNf14FMX4Txni1XY+p0zvshEj4b2Te2Qour
4om6/xMrb3ADIZxBCHXg5pYYhZmC08UqjuTSey5NDDlHNuMQMwFbkJuN/JS+vt8aMXbyNb2ga+XL
Oeh+hJOP6kphbdXV7pIeXWBr8kkPv4ZMrpcg7qCahy8bOklIzhWderUyEu1T8RlEqU1GQxDTWaer
aNeMCrgDBRG3qRjxmC1b9lOiGZ37iGVlBg7qLh2Ddj+J02GAMLXm7JaCf8aaeTBysg1aT0YkH4rB
nl4jdxsYyKM3vspdp4ynTdubVCMhBiPUaIEOZ3EF1t14LvOY/cb8DRepUqmFiZjVbei0X486ig4i
QBFuHSBSzvPQIwT0sYIUrODjr73be2bECcsqdkeowar7mpXn8jq5HpyUuiHKCC03zXB2Ut9fJVyC
h8vcSKlzcOaPoCqp0f8CF0faIDhB4mLcsPYYngwpGhrh/VxIcjCACbWxAmIAiVNj2t4AdtHLvP9t
OvXlHVWRpWfEuCnx6Js3EKw9YvqfdyO1+KPuib5+4G/1iafHTyfHGsKG8P/+aiWwrvDojHUHZh6v
rqPaLvhaWJ9BBOcEN1F5LViKXoNifrJd2Q7RNNfPuLOJpOUtgTxbJx1SWNd6brCDfz8MIwTNprbt
MqLOui1+oQXzNHPzBAKzT0O8jcOSJfNG5xo2fMtCVI+wE1hMoUvZcxitbP7LibprJBzvXdoZqz3m
+prl8vGSeTNItwtGMctKnjbS0UaQU7SxLLtpmyxo15zFfMNqG5VTohEHlsNxiyRsxYHdihDnQ1MW
SGT8g9ReWZGEzsLTLJu0PeN2DAl3+3sPvjhMG0edu4wFeYBag+qWN4tBkpI3Dcu0b98V7gOb9iYC
yiMllN6naksBi8L5YxTGC+z81UpA3TSHMHDEgJuYYb6Z1e1d7u5h5X9nnzLjy5BqjzKFaJCzF1rn
MpvKeC4jNWSCQMbE0X70ejvyMOH54Ki9cASlvICYgD7XR9A2jZGHjtMoyXa+PG49+9X9/6xjQWwu
2Otq9lH7ZIHvshNt6ChtcX22Wy4xSZVhL4u/0851/tT8nItZZcLiah8p5Fr3JJky7GQnn3PePKn0
OS6AhKnFJ22yGJAp+B5rnPBblHQ9IQ6fO1x+eTkVnJDjegiaqlEDMtDbRW+5+OslLpvDQJEFIk+C
7MTAgOrid/cHz3upA/JT1tH7+QhZPi4pVHiZCLujllovq7VJkIJSTNGl/FLlq9Vg0K6116zEgp8r
dXGtrOXASmUyRoO1Ar87P7DSXpGHhHm++e0b1+/9BcUdLC+xW3EQs+8780dPdexPmt7icxWTHINq
iCCyToir1PRAMPYz6DD5bLqlQi2mqnnrhXu4Cei5fIkJTquu9QJObFz/576hCsJBDOSBR3T5fvCB
7dy6E/VuCIG2hWxEf13Lii2zr5nHVVLlQ2GU3U2r76Fd4W6GL4655ryZL3f9ZZmCXz0T9Z8Yx1Oy
y2s9rVNMMRyH0OWmNwI06guKtHOwf2U4UBcnezkGUJC0OOIG/FG7mkKdzbVOMu4QtmtQzT4lbHiL
nAqrn8VZp9U0mH7RnwbXcQb9CdZ/vtHxDP2tmYhJrGm8wOAhGjkTK6f6GTusC1rze/nO6399h584
weoma2Ik7Kbe14sE9vKIzXNy//c/jVjRlvUnktmKGcpBFdMWRarG+V8c8RnXNK1PnwLO8kn7LC/4
OIHaR7+8d0lUTHuBZFrAaeGIiP1HevAhmA1MHmbNpE2cufmsTnb7+2hT7BSLpUCkxZxN+TAUWofv
dK0PpcwmG1e9YJF5JQapKLtPWelWKHiBoqT0qTrdD3eSTHVK8IPW7yQGhuP19T4ECKe7ebpchkqV
6PDApeEqF3W3p5RcQ0xOPLCZkJny+XoVZRWW50RmaNFEDNnqtjEOS5J4iQGPA5CFmw54cwg39g3I
qz17M0plypYcFWKHhAXAJgeeayChw3Xn7a8LE1rT5TU3go2Q8MUNChdNbhsQ6ULpspMFyQhvZhd+
rgkctiUKrYzvJOxy0l5HCXlGJ+q7QDfcTpum7mvTPeDq2+YUTr97CE8Ey0iU1NxudHBXCyiNDhlZ
+oVkjmoSpMHleH0syhCWca6HAKOkAze/+uHGDD/kpfdmehPePPrT1uCKRt79O5C2aYK04sUd2PlK
fhVe4iMr2ixluRlrvNkqLE6w4X5gkDE77fAG8wOHbD21hkt4htlf3a/vHDs50Rhxm46x0b83xEBo
1KT6vL0A35YJ/DmYRn/rxWvNrIy8AoZzKsMdWd1rFaq2ItH9yrWRhGJNViNoh5AjnMrkX7thun6V
2Fr6A5VrGbuJRcUnnx4TWSnewfQslUeGZW7ipTtufRekSCjsMkgvLkj6fWWqbaikZHen9Qr+HfK+
fr99wkZ4INJ1gfpdixGBKe86Sk+PWezKZlYqPO2dwkiXFXcPcwF8eG2E7Mw1sWExaulOTwOC7HAv
nUspxCaN0AfWhY5n4FGvciDB6cS20ld9SyORxJOam900EVWaUFBr23xn6hcgFw/n09kR6HXlmHsu
SM0LnmMNbsAqPgKZQah0xtnPkR20o7EVRA8iTT5CA/wd2f/cErMXb4Z16sd8PRaUgJfjyF2rgXWb
fRh1VOC85EKAXIYyM2MX5zyPTJazcgfH1phKxf4YbSrQS2KGd+57NAmnIHDhWBOF7eQPT3C/Fb8Y
jBKf6CPjT2p05L+WY2DYOdB67DnPKDevF/JCurmlqeCXNwCIHhJDS2cw6uy5HnRceNkAqKPUJXFO
ziyxVJ5dN1vV8jSnZuiRQJTeXWQAV9dmnKKg7/mjg/2H9mnAVmmfiacHJwnZUqin9dkxwJgR3Jym
M8wUxGanCZbQf86Is/6DMAG30O4jFY9gvGOGIHsW2BohzwF2C+OXu+91VmLAqNYv7vDjSsSiRRQo
e3g0VX4D8FRlznkZoMt6cEMA0tvWiTj6eg+8WrRVvlK7bukUtJkdZEhk8PpYdnrr96s6JRCMpiRh
1s6A4CVutIm5wx1FG//UwH916TKWrnW7xa+pVXaeLB3q06J/hG7DN7TixrTNKuPzlBH6H08HyWfz
ssrw/ISB3HQnsvIYyj86mDAMgQQn1oggM2S+dR0oXldqzQxSQ1dhKLx6EXNBnlqLZRvvPveyMbLf
RMUeRGq8AcIhn+VjeCQmYIjkr9JjXe5A3sfpGFkBgtziPjTk8xBTHgqq3ENXzl4L04abahvenbEa
EmNqWNsgXl5LRHfLWYS1Ie+h+K3NjGZ+Cy2slaZNFqyfNg8CYdKxel89oUPBeDORy6ifHz39S5NS
ipjLHuThNyJvhamP1H+u3mNtO0PevdoVsCF9wT+pZZaFNnb6dZtjTXFHnAMyw/W3die5mpNQik9y
m21aPOmd3/MYGu0QUVtkhhU3GvZFOmdJWrX/uiGEmuth4bdgmsHMGMcVcidn3H4S1oVGNmr+O7/r
RvYmuCCJQ0tG6iL7VOqwqSuyT1m/Wwhpkej+hgJnKf4Bi6Tr/LqfQqXnc7YbW0jDIBhMV7YpE8tm
RvSBtzaV+HznzUfXuWMqN3skWAmoU8NnZAq8p7C9h4c0tXR0K/nM2l8YLhKG4rlVGGG9S4Fqwf5C
ujgkx1wDTzyq/jfv34BP0zxe56r6kv3ctg/nuitQ0RW7D2HOpubK6ysgmSDmluCFD6wZpsGgnh2l
TqNr2pdyEGNZ7v35+/Me7j6EMsrVLo6tMEOV3PKjSLOUKDMK+YSrJEGwDRXfAyS703DhG2ImCjRv
wCOUZus6LR0b+nJa3QfZLDMeZ2nA6UU4GAHXRm0mO1LW4WMTFGIx+MfvLyK4A4ggL9sG9Wre4deb
tXYkafiSHFSNbKEH76qQaHV23jCNc5hKU54buVrSv7Hyl9qGyzz7iUlH81Lv2XfxvoK5BIngWQeK
dM0UiTMy3dI8vpyWGBDVxNZpQPnpFG9VggI4pYq1OFgNZ0qn8VC9Tw4mjLUS0+8JNwvA7/71+6pn
P3EZ7HVVDmQqEwC0LXUxUUc6XxKcJ/yE3krlIxY1TRdUIjfpy7waSQrYM5O/7T+IAFRH7R15ipjq
CzaZ0QVOElTqnPuihX3q1cTH58JGXeJHjm3AwSqakz0Wdc4OqzsB53En04iOh3dIL8nfm0UACUVM
7rwjnUi6TAptpsn+Bw3jOeBgk8XLiTsHZG3B002yWLerVtJM2gaDBP/hsbvKqOubZhDZyZObqWzg
gw15FcOhhVuXebLSfn+29IWc9tOBV+PlyuObs2ykhIqynKhM+PWUJuIU8k2TaV5SdNnQOlF4W6aI
Yh2bVUxn2gNsM0RiZ/1RSO40X7vDup/Rfxud087qhWKPITPrtX+EwEOugo9bjm4iyVX2ARIAHvqc
27PqIAWt5kB154MD9MJTt49oHXJLGt/ST4zm9NO0UX7kWFds6Bt4bFvchVxzUtaxqBKUNcBiTYRf
LLK38MTPWzUQ9qguoeQCAHNeEHvCeVQC4QzahUZGKgJ0yNTwsPa81vgUfBuReQVkCzgbTS5Vg44s
wKQPnRjOcL155OvIE2dTgv+mgzzwQ8BV5Ahi40ujrjDRBuQDdlBYlQEtoDB8vXEGnTNPKiQyaw2z
J1MK7uG9EHjGmKEYJ0Zmdrtf4LE89lIysjA4kduYM8xBMOE7NcRZ7PnN0Wqt7gO0vBIffqXORd62
YIIK7g1KCjRiEqqVyTSwYESZziqTgQTAjKqarpYk1CImU5K4SyRKvLXxbQCHzy/Um5+Y2/Kw0IAX
ELGg3j3eE5Gq9qKaRTKhvhsuyST+dB3yrLPcaaKl1/SbygSC5szQzFNNGHMgJ7uMPEKViyIUkE48
9/XTVdqki2jEiEPXBI+BE3BHxHQpz8k3+EkEvmLpurYp4bYWSo1/Qv1HA0ABP6RmOLZzaRvQDdAi
S+9QLGDX8FQ6lBdKzRsq+CAfg7Dz1JxP4X+9AsZqBreUJs1AjlzP/k7vgsmwQEnVxBfnvPPyXfjE
HTD8qch0gyfq38I/U/oZvsN3CgajJPbkmWZrysBG7Gnx4hwmH4qQwJSxLPNoqVmPPgGbyBebnDEc
7DhUVl8Fz40Kc+1CvgoHID+k+x7EEww/kc+oATVzGea3W5Eb64i/KD1S8+F6fbf00dukeevhaxBc
S32ojp4tGnYDiByY5pq+iIdyhf8djOTp9ZTZV9l3P8eMbmH5mm6ue+NzSbRmtqCeHfkx1ZaUS0Tq
dLLAZyTj0gS1kQ7ZQaFyV3baK382O9RsY8iJ27ApVQ1lBN7WUAinglOviJZssp/qr4TKhrlLLulp
+5LimPYOkURySfnv0vYMZtMw2zhNYLOLjZA/gRygVg52qhJ3iwgNTWczHB671XyYrZE4u3ykCEPn
5s5qagW1O1//OkmSib1p/sZ41KomObeCdM1Q+Wp63dkXj/HCa/zAKJeVPhMopGx5QUTbNdrHkjPQ
YAjQwW5aWCgOtleDXOfdAmy+jR9g4bA06AwCE50c1Z0dz8DoIxpL2GtBGAfu4I8BcNt2QQ4jq3K1
xRCqRLxy0N78BFqFDuxKdF72WEk3QDmHJg6igpYyM9a/aydTCt0v/Wuj2c9auuEr5rETHHjnp1tr
Exa5yTet3fnPy15gHwJT1HtBoaYvEAs6EpkPb5CX+jQDiClQo+qdKPbyylHrLa7cVBpZgLF2swg6
pugpwJ1JuoSJcrlfLx11X/yWxblOzGbwcmYLH3WS53uX6/jDEtRhfpunjZHpsY8p9ETpkz5WR5Cc
OyhJTZ9yAITfqMjhk1X4ubLpMnK+rGA86a9YBDYhTphul0vfZ3Ocagbjv1OqOuk5mbuy1Ww9uUX+
TmPXgEJBTyZvnuWIFnRXyjCUgKqwLWH+S8vd12immsPA2UFA/AcN/YxlGEo684cyk6gaw9VAoFIk
MzNF24stWDzAPhgMyw7nMozmEx7g8uN/rYp8dJ+pK/EZ5XiCWu+uDHWKRQHC9Ys1dU6BOBOijGKx
RqVUgkIL2Pi0xsQRJIWbDdynQL++kh+MQLyJMX8HNof00Iosw2Eo7JhdjTuAlPLeWTwWWwgNjJNa
uwIZjPqeTNyaoawLzGbNdbVbVxFDr2ly0fqC6ZmCo8fFI0vOi+fi98UR/6jJ+EKnBNsDx7HQmV5N
OJxeJvgsYC+UODChXLxvSsKyVjDu2RqDekkjoGhGaanJHz3WCETt1kBQ6qtVQPo7tpwhTd8fll4H
3LFvsHxNnKQUMQZg1eNa/81fD+g/0OANTVIgw1QaHJpQ94n7+jmxJw5qjbCm9enLrfzTOKBdohNH
v1B2jfxugN9M/v+Q0oEFcZR+R+t2egGrLlxuixxF9BXj0xxmV7z1p+tk5y3Gb67opKIgTWHp72dx
feRaeH50NWzFsN668RKZ2VhU7m0lCf2D
`protect end_protected
