`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
k6ZfVwSszzfVs9nDC05c1G38lDgdIb8KnhMryD39IDhUg/cXJFxM219cacsw7N2N0gQoiQgEb5Jt
U1YFycx4Kg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
M3E2Ywi91iWZ39T+a52wOHF68yAhqLJ9BY40dsbNA8m8iWG8JwUvhY/xmDdw3UNePQac5HyYrrr7
61AwwRsfcYSkKkEEPeCc0IppQArCUVWu/EPgBxMKzk2vEkcvibjq8NSWSpWlIq+guK+qXNOBOMOA
6h86C+PD3lxM6hkMm00=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yDsULOzCBoCFO+YinwFUWaJwLEyD5/inOj517RdZpb5tODEot36JQj0771r3SFmNki6FVWDhYVG/
OHjkREfyl/ctmgR8l4ptXEBihvcHPuliWqtnw6lCYGWwz+ItrabYS8tQwdUAYj+VyHHuQFUgAHG0
YYASPxD+rkNTkGJA1Cs=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hTtbCUl/7TITxb+Dg5Dj4Olwx6hg+MMuhtLXdHsDxE6wvrwhLUGNRdJrFz8H4HqtPuGYlFn6NPmX
Zgpic6yd6sP77+FGnGmGMBWVOLj657vecbuHCrVZpmZvIiiWPXm67FLll8AxJZVXis18WHCo2lJD
5FlYtGd33+QsFnPyNAxSg4hIIgfYhYz137TdcNQGCQ8N9vcX7nE63BAdgYH0ol9LGm18OhEKWDOE
0b256jry1oJqFTf+yc7abz6Zw3wOaYW8lXOUhpGFBOY3olBjkIN6UnzcxEK1Iwfi0VQ/Tp48d+NM
w2A3/gvNTzWFAul8pzdtqFcho+vs3l1j+4sL4w==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mNQY2wwnhYH056U6LW3sE580T32Jyo5U7MLrzHcvRD5/pfa2RjXixvv2G+Os6XySDSZJvVGR+Rva
x17IVjV9v5QIYkMvWw0NUg79UuozVpcmvnEMwWdHXixmbgUewXlQWq8/s6BNEB3fkAv/W0noV2dr
fJFP5BLGAuO9G2FHTdLHStiJEkFTOglMNIjvnAM8FSYMQK48uLM2jOea+kC+gG+rdZ87sKvgUeQz
j3tr9GRF2dFzNyF8Gx+ZN7VmNur8Rr2DWXcTMTUgkg2/gqCu3pjVVCOnLnYt++hCQ3DFkJdHzN7v
NeLqzHjWo52X6kbB0gddMo0alcguHpKb7EC/eQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CuhN4i3iT0Z4GDwLURTtEJ0A0kXw6MKHOkx2V202b7PrTZi9DYH4Vxke/sKvwCtWBG7xgOFdsV8c
8+pCSQkbGpUnyjRtvLMbHexyuauu/DO4lZYzZhNYDnPRTZZh7FRMeatou0HOpciy2vv6OWc6xWd8
SwAMB23grqGrnML1WUDOnyExASwAPc7kIJBZA7MCpNhJLpC3Rv5fBG2spHqTBB2MbG8yrRiKRTQb
huQrSbjsxY0V0yFBHZGoZzXU+3Qq1nul1s5eBSj7kYq2jTAHTpacBHK4JylVtg1MMPK/2PyTHrl+
HdF6H3v24JzBo06ViW4ILzkYhDaxmsDHlG/Irg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 648640)
`protect data_block
mZM936nOMJaiFUjeuBdH0rUe7bhrALdtXJBn7eBMqQeuq9VBN1VLsOyQ5F8cqvW1NLT8Uhw2xBGV
RDyA/gKHmDw87j5rYgaorOWp9dAe/whsxeGvQOe3Qz5sY17jFVg0RFFuIhFsnw8JgyFZZ2oqcbM1
AAvSsAKwMFOQlxt5cqNF49XhmV8yCcBkB0Vbzk3jv1gTG8ES6Q2MrF3HZWq82eXYlNtZXtstWRMn
eMUpPUyzXImdBUgd/bvPWlaOURm/BAuf6M648Ipe1u7Nnv5U+y3ir8wHtqyrtEkjiLBMZvT+a0YF
qgJatn0CbCxSRStbp65o9WHLonTXD1XlFoJr9bWvCK4WsvGVzyVmFpKwtOzR3H5NgMww5Kzyiivp
34wW7Zb4PvnEhBU92w/kVqnph18GSxyqmadSxW54SV0R4vZHXTXplKlx18IDPqdhJrSz2fB8y/5V
rwLA9F4QQiN44+x+jwX67DAyW6KjHlXyOFZ7Jvl6jsgI4YQttXp/eW2Xco2JnTGOLYqkrgWNeeMS
y6vsSzJujOMTmP9Z3K7NB21pfWxGkOyB5SYCa8Gm9g4LiTKwvWs5FFg+DkG3ZAJk/csL3D/uww5L
+yrJXiS8vFyYbK9aYNMI/acv1SL7kMDdhFzCbc0Sd0WEDOJ4ANhZphSqfGQ0yvxW0VjJwUsmmIXO
zOTixCOIopWCUtN+NbI/cj9ISCxcSZS+xSXrFSMQWNnAouEfmo9rRgfQCoBGcIf1s5hLB+cN82nP
d2nAFGqyGsePvo0VrSofSlFvsdoiRcuZXsYUODA3vLcgqzVPuEqL3wLPfbG6F3P3CdfWz6RF8/Tu
IfsTMMwpy59bRz6CBRj2IWe7+Cv9PiGCuAGy07E4UbI5kJRQ+Atyw8oO/vynr4CD/X0aucAMzNEG
7KDbASBFVeLfU00d6Hk5SUfslP/a7GZJsNJjBV1CbQY+1B8RJ/jYBSEz4if3sQ6WIjg+afstzrJW
MOoZbrrZXk8OU/r5Xg1bvBFjqaERRp4ov+Yt1stF6Q69QJlPTfUdGIWT6x1iLGPmCKBDigYp8dXV
S9a8yQbUc6MCH69R0k/Q5ZV+zkzulXbRqPszYbHLjxonv5a1Nw7j65+nEi+J5/JJB5/qglhzWqQC
01OUSi7s/h4kZJ8sCTlZEfjpa2WaE4TUboggP75HrGNMZL5metAFUEzuhh3GBu1Trrj2ajFlRcWN
Hsn0QxMiu14lOAODucYxMlRMzTpHGJKEh9Dg1l6UX8zFfLACp4vVaLWCWZrPpeQGMuO9VguEmvf6
98apok//sBBQmJaNdxOi/MF3+LI02pHBI53ysI17YuQOOwP0uohmyny9r+n7deYK2Yvoj9DIp8d0
WgX7NZ+SiLnk2CIX6XBDubCQOkOJtXzFKzcMSCa7qb0WAaXH/qrF9K9I4vsjYwPUzBj1jqP/flCi
+8x7p60zXDy9BT3YWJqIWYOERcE8x7Qei+TnKZaOwxe2a8xH9iDn3PnjGVvLKsxIMzGkIgGxDLl5
HvyNFD0rlKZSHf150PgYDygQsR/N7zfh8R6ZNDSwRCiKxWAGposS4eRLWTF2MxOwaZwyABV096v/
qlCMXzPEWALgcjztN+WncnZekPvsB985kboddiX2/o0uYbhvH0r8dLBmpL2CvHjo9UMr/TkJAfjo
yNGZrIAxF0JCYZnqNGqejoe9gx5wtG6ag9jYWzB5qBMl7eWRnOC4Kx85ZZIZcjOrmVBk3Iu+Fn95
zK9ZkIwuMKUQGLJyRjLxKUXM5Po8DKFjIz41GXsO0fCN6XMGHpOtj6WD9wSUibV6YhrUOZCLbLrM
uYQn+ZE4VVqXUZKTOSH+RlrQFWPbeKB3IlGznEpGuu1RxDE+Gzk3C+vuGpZumYrYuElNsYK9Zt7L
DU4PdwvCmrChAUBEPGUVtgMK1LSR6eA5UI1nXnLTvfUPRbq4lyaWYgkwkvk8EW0RJ5Ff/hzxnrom
pfV/hnXJ26EjK1t0JiUHQtmjWG2s3usG5m1LwffTXp2WMemYp6T4K7SRcMdJkwymj7vTnc1XAkfO
rl8fcp0FSWgSOEyVBuDTsTLt+aJfZZhynk+ZzF4JaPgvH4Tc6kNuaQVinIFvomwFJJOMAR4mYtd6
2heYR/Jzf3KDCJH3ijzy3XsYelU4jJrqRWLH3N52qQkssYoLF2ZFRCzducOEXzAtHfA4cHCa4FY6
LwcOKWV7gD7ZDhgQZ3EVg/7ECpLkUGe2J7bp4a0cwjLQ0mMjuGditwIksmBffnOBCcBTZG1ErIM/
uGL+yp5ulOV0EmD2XL/XJxvANR/jn5Zp3/qO+GBkjeFhc+zUuq4YcTtpsh2GSHDp+JtIGgjwmjmh
zQc7IhFabfmqH6YiXvgo5rgjsuM7VUlrNsGpEu0EHsyRipl540SrfwaNpD/m2UdThNYIouBwJyLr
QfproINvxGl/6g2jvBgQ4k2yF50fuZ4F3O2Ti+dw1mrpJIjJ4Fye93I2HrXM8t8Kobqff4uuEgKg
Vg0tgt+BpWDEy2knl++z9vjrvsbvx5WxPDfmWkX6H/IudKv8wIjIv4PffUC7+o95Dd5u2yOuBfkz
vDTu07ONVJ0AIYIo2dW0Qq6sOB5hP/3C7DBt/6GypB+piCM/A9zAhLjFG4BbZMC2o3xV74Mtz+Ek
kZvP1+8TXssBXJHVWKWGk0JyIIwZYkUVCpSWcARuCjxEt+rjRV7E7K3i+DfmAa//HN+B6hQfMfZw
Ostrsqgzzgndv3F2tKIaeoiGLyB3qYOMRuCoQBG5kSSqYZwWTRT10wCgLOYlx5vzH1/iFheuQjAV
t3yTE8qVhZf60J/x/tSo0HAQbEWtFeGarQ4uUix+L89TeuejhDGXIO5lmWrMCrJ9K6+5uAmTYcrg
4/CqHrTL7YvtGJL39vyOSVe52K9TvD1SLFXx7ojSimiNjCXgjxkr3v2hGRng4gOrQonCrIm3kFSF
DqY+0VXGdlYfLz71kxqrxLAoHI+74teYgiAoGckVfjQSYNA9Ws90xpEkt0tlBE1ri3w1rmsFYdZa
yW+Ixc65NmIluL9FyJBLloo3NNzCnvZL3mpsn9IvaMTWJe9F0X6b7zJF5tLzmxsj63Uqo+qJJqSu
Q8jkHC7zGRWGaf/gjnoPk3r3VQhgKXF1cMpeVYZqhiT8HGU8qvG7sbpBBtjRgzKGzPfjp5bBVuD/
Qye/B7aU9d2OTexOufDKY7p6WMs/tv21F4rzmw2qQ6rcAWa309Uy1+dFwJ41Ts28m05/0lKnG7Sx
UdYuVK3NVJP6to2KbuKP6QkZJGzq7xpQFqXdUm0PiGlrovLnYWwDayKVsW0zHsABtOFvpl3GAMcG
R3QdKypoUJl0c4pa80K1kx/9j5fa3hrfGwoVTItkQSCPSo1ELMsyyquuqdPwwVtVYGJThaJ0PFLR
px9H6UBW7jeUK+m9iCC7R4vlFWUoVLBzcOvO+fKkj9s2LC7ENhi/fhycb0gdp90ztzXUZ2cHjqhL
uTfNvWM0SYFs0I/Lki69o/TLibfxYZXMeuYMNj3Vbl+0Iay1OVfV0Foqr4tE87YkRF0/j1BhcuYd
E11YeuEj1RDR+WHAspj1gz9oodIl1kO3D0i8kIlPfQyrl1yPD8XTsr+vPdOZIndlq0+qHipL0sEG
x1na7cgQKAKH8ShJvrX2HY2zdCp0hGQcFmnoEpzrcrENb7ZW4OQ2405T/51b8azEw5+0bb+YMHqD
rVwz5Iern0dqZlri3e7Hr/Z52PAA4YtMrdPaGhuUgq1zGuJqcySNZzTroV2SDPSdnO9cnQ+MTfjc
CqOHpXbyAWjasxpGYBw8NmHKEMVuZw2u0XufjPUnRLYF1leJ1hirUDEXoeJ4OQzMwOTQpPwOv6Uo
10oMd+aGsn+JLAEMxV9NgmH758U/0R1aq+RyQD3gPJuO7yC79csyiCaheYXlHXElXSwYM6dg/ozh
I4Y3m3kJP6ZdnBcwC8KO4bWq2hy6BaBI3sJEqKsCTsD+H8+6ctH7PlSvXFLyBaQ0UFhG/a/Ajy3E
xXMF+a1HDDzPrcE2LHw9v+h7W628ocS6HHsfcgFHjS2tiQQAlvFHfFYQ92EZ5PjUlE3jdW9jADOi
fo9lzpSzwDeaxM+q7njh0zHTH10vDJmtM621m26SMuEKfhdPg2ma67I0icsmGknk6PcoVeD2bENQ
mPCiygbNKWeqmovSsDo7GidWfuyzRzAcBkqlj8Xq9dI4hEEWDKbwHLZ4yq28JaAD/J+VOZAOWVqr
MNAh1gopRZr4P+UifJqSFSeo8qriRwMbT8h9hN9yE8qdf3fx0AelYZ11g4i1Q1aLctyN4m8Uiddq
QrRmQU26b2vIrvalPN3QxT1sQOoNd38w71Y7e3/XNzyFLG69jnBvhASNm8AAggjr644HSHxsckD4
iKrV0SLcQ7g3hhNe3s+qSJSaWSftZXc8mWCW2WTkx7YBTdMjzE9w1VLori+YOegZ/Onba6Rst5PU
rT0w83j3C91v8cichnfxn5Ga0Br2lJ6h4+gsRNX3Cu+vCyNfumHDorGHrfSE30i7gIsCo/j2JRB2
lr1X2Xm+RXQVRpDaPJVW7ol6Arq43uvj/b+h/1b+CttDI8cRC98NulxYUWDtbTC/v+AqhgKKpnjV
Cr1Nt90wkxhHEcRndRgSlbYmI5Cue2sv3RjrXRjTCUeA25w5ppJE9xZbIc3DOF9GJyrNs3GHctZQ
ooTyvozSWU3kpiQYlL4eQcEvoti8one/vbZq3vgkEtEIGqGv6wIBE69oy8/LHGwKPzuG7nhu9+v3
vpXRO6XXAJycXPMxsP+jDXFmnBmhARfUiK/4m9xfjYMdSGA2lIBI1Fs0zhy0uuwDig/NDMlbcRX0
oAZCzge5vSvE68PlNJl/YNUK5VjevrzijF4+vMQFor8oT9LqYZEoel7besAT8acZz0EahSQi4wqS
ezXi9ZnfL0Fa/hIzI9ZxAfA7aWscWxBhpvh2btN+37Pzx8zn1RofvS6RewuUj6jSbF2XS6qDrE4y
aR1WKz2JkpJfCmNHxYBBb4gBk3W9pxVScYi1nVkBELmf1t3wiGhYyEwzEuovv7JGB1mWsWDuUNFW
8jrenz6a7ZrmuWyfoGkD5lpsKjHtF8Iw9hI3SP1awYjlIROzfTAyuzbt0uU/7Z0517ZtigJxNqOL
6oMTX7kqDTvjc/g2sBTwxICP25+xYYmrKLE4taE8PRzFyTTg4dpvOI9kUPzs5IioxWR0MZIM92kX
f9FXrcFjYoXTt5FNUcb+X5RBUuVUW5sYGReBd2eWeVIThiTtLE1Ekz32y3+tkZKwTV5w8dkA1urA
eclXsRJ7oOLsl59up1HEBBk2/6THErr+1EGw230VwzP0HCPJF9E2fvfwoqgRq9l0XYsWmqYD7+wC
ed4VlS9icNT6y0S7/aN0RGEEpm81hOWou8zMcbzQIcn1wvBQcA7K1MuI7Zm41fPc+b6OxUEDv5aL
o4zK+PIfKFsYimdc5ud5vULuw8qsLpkRJaVHqFJCKJERSSs/6dazRcsr/uPjZJTOj2skfpsqUuxw
ugc26aq3LE/eJF1h7qrIOMwy8ygigVwEmgbDi/h+Co3oHOdwtqGQh24/CPrFbRAfy7fW5M7CDZFf
yIx3RyzqHpU7zYh4XY2jBoRnDVS+nW+DOiU4DO2zC42PZtjG+aZmFWPQnCOZ6atWoy24xmdeccNZ
9Z5vIt0+zax29k0cNsO1uUxDz7JJfFA9zTy67vWnVFqLZrpM/ArcPtTOtV1guDpCks1HBcrW36AW
dCJ9yaMQ5XBxiv/NZNDk3xAp77+CCeQL3Ax2/toWfMQmT8Is8V60bzOW5rbkMyaSo4WImQxokjl/
HAjd5PtpNRj9NPBTudAgqgR0UVjq5jdCv5PsgYRappsleP6KN1XmuD/iF0Mwowl0p9gZAGOU7Kl+
hZCsOOti8aMwFp6t4kKMnOfsFmomygIpOxfYVW9BhOsnev8Fvxos8IrhP+8GgykXOe8i8JzgCKum
rIbaOdz/a3lJqmXkeeSqwRxeDXkqaF9XbmLGEmpL1F+O6FJDdpH2b/RUMRHiq0Oi69LSMgKzauzl
tcO+VAsBGYTAdkLvz/rIMuyKE1XCaCSWWVPEQfd47kK1vQleEA3ipjNAG/XJWiUrMAEC/2Sp3Cud
dbQtYI4F1od3bR6r5tWhKfqemwHogpZkVaNh8OyF3iaVrztX9b/B7yiSkx3kiz97JcnS2mdqDk8D
yq++EuJkiiyH6r9WTKM6/flfjyTWchlV3Vzk0rNBMjngXh13L94wlwpmPZ1Twyf9V90C+TJW8dqu
J1Ef5aWwBIexfNGI35I315+RiSOCfDKnHISD3x+5RGwqEq8eVHMnWXR2Quph4o2aauMBCrUfFZG8
lgdDqQ4kaNVkYvYx2TmfFZeoqmw0+zy9fNkMGaL5yaiMaFXYT6YurOdxfIeSj9i0QEuFwoYuMyBE
0ESpCdRc/uduTDKRg0COwlHv6RbcpUjHurdFChKiuZ2/EIK2kvnwlOk6u/o8cNqbnJ4CvXz8ZbKI
DeOERR43PwQJrQmvqYIDQdHYATrVzFrEQs6pvhnvtP5mF2sTm6MmBqB5v3J0kac21GiHCe+nEpj/
qkw2pq6WWKOdAf/mEH1LhPkEf1V+G5iZbZuGbFBme5FLs2fv4lBaRsGK21faN7tAONxKbY4w9slN
fv+VSNrEbJPHCwAxGPD6fgG6ar26+dsW+Qi7Agdj06gD7iPgTYmDCBOEDDp33SyaqSBtjhZfe+Oz
vCWgn8cZX5JAT9ANL62LbbyAfoUFJPsPHUqfSdZO57txgSUMOD7GTNh9vDf5xlRdb5sh1sdWDqZc
NXKejSoJ0y+wqsGZC7NLc75AOpkGt0nrM98dmg4j0Eezue9yOZ5DiB53ioVv2KccKMPDmzOQbokH
rlgkyybwWo7mL6NauTUscx9WMpDq+WPHsrfb6S3mDn8eiJAvR16jvb0guoJpIJm+qq2dxm0rKbRu
BV1tcZ6nbZVXS+EK6fcKw3vsEF+SFCNI5YPLNA4UgCL73FXpJxJkTnx5E2Bq/HEPIvjWZpYMF2Nn
FM4FC8Nj93g6R8atLqw/2olxNqncB+UOKLGzFa+4rpas6/KJZsNYcNpiCDzTrANh/m8BKgPexIsj
BVCIDr6oDOy+Iiz9GHnYpm2LDGAgJcCaxOdoq0RtaMZLEr/jJjCvrB8wesZj5R+AdLV+yT3Cjw4F
6Bnmq0G2XYQUz2V30QpbyLB1q3PNJ7C+nHeP08J1gHAEJQ7bHnPuxjl1bf1TKCi90XmOv7D16NWL
244kYRF0VM9L9mNKKBsFPDK/PB2bAlOvsOPB/9odqt0aeDbBLWoC8TMY9065Fwj7K9ePqOaeQylm
l2ZQjDFPMHznP/LV+UWncz1UfmAarhT1hUp7VxPZJuV/zTZ4FFBs+h5PNmTPawm+ZNsvg263RSqL
kjsh52LeT3qrxnOU4hPEdTOx3Ll4XZXSnf8WrWEGYig7NdiIpZWUhOOhmkwp6BxStugEKylrOlJ1
mxUmytshE0QenD10bgJiwiS+2uT0JEV+X1qJCSjBTbPqh1Znad7E/HBhRKBuNlkfTB2bZmSWnWHA
4Rhvs0i6Duuf/dLGBGGkY2LtaDXVRswYhQOMQhJa65BlROl16UPXFQptNzvZSatTmWeHwKdOaIgm
zDu67TMPCBnaV4rnk4Jz3gSEyzHoIRq3kyuo2Un3DNNivZyI03XTie4hQS0r5JQy1dmaWrpEpzuS
/wXYL6DvsiSdroCMCK+eakeY/JGMYkda0zlflcJr/1pEUoeuiE/j2JAc9AYf6HKOsIlaPD4R+Jtq
N8+s4sxI7NM/nHNalxIsjSGNAyOs5kxKGVfexJ4SbPT89N3nHktXQS406V8w5n2F92htECJu4oU0
aNwisboNESF3fNt2eVz26CZu050OtfLNNMK3cFinM8MBogIgJAubu4iEt/eatWPydhfBrb0vQsp5
yGI3/ZU+J4YhAnGIX9qv/hkokmlVibDs3npwa6l4eOSXSvv2htcVI3JDbRmP72Mw9FKhL/oElzla
rr2p0wa/XvW/LuoqhfEcrH9qfxIcobfqNw96rJONR4ELYH7ZuR5rW/5a1dI2dTeXt7zaPTZsytAZ
wuS3OCTi/P/kCVBCjV4yBD3vVhD/ZTS0dtQ+aGUtzOsegrS3MQ1Ju9pse+jP57sIpPNdTB0d3TWr
qOC2253T7R/bZGHbqMy/sJ5UNLb2+TzVkQcWgumCqZ0JjclZ0g4EDvzIaDM61s6WVj23w5LG2VA3
sYgtFkg5901xjq9ukR4tAAPeu5n/eZw0lT/OU7japCoMv3a0PACXS0xRyhZjCuyEJWPxfPE9ceoq
3BQknwEoOCKNmMA4bNVkqVUO6xgFIeN32C5DYH7W0+NDqeMFEK8UgyvO8ZjlclKSaQ2nvdMU4xnu
t1m2ijNnoouU1ljatgCucUN59CtLlThgLloOzuate49Jvgaa7WzCWfZmLy6srmMIRbSKraQuK3cU
PKSSFWdNg6UN9RSJCicrSy4YJIdxd7XzQei7vn+1gkL5z1d0xs6SLBcB9WASw0jfFi4/lFRzmuiO
/ds3TCWZb9Gp6dibFPR/52bFeBi4SqKr2XbRbAuBo3lxBvEwGtK4+dROMoKeY59zGTDGNvC1Rc9v
ExC7qF3FbqYsasYGsAaLY68CLl4j7FJMNqL5cTzlhM2BvdCx8MstZxAVrww0Y1xZtgqm2hRRSksc
8jRBzVpo92BInSHOoJt0xbGvZqEu7xdpmURJ6/Abub26lJ++iOHxV0Q/UKhDy8yI84Q0xVjx2pkt
E+s20y6USe/t7FUfj5ABweX1GzvjABEQd0AfKpE2z+s8bRLwFYx4rTvLt8287AA1jkvleAwF1Fn5
xjF3zy8Qivw0YO2OXFh15Nq5TBWHuFD9cFOzVmz5hiOfrOAm29eIIECE4MqeFTf4GtVq4drUhnDb
v+WKT7k6S0oDe1yd4mvSV6RLIuvm4NtQ9Vnzgg8aLruaSKc6HM93xD4BUSmcmaeOhalhu9PDWLBm
2ETC33NsDIGf5yCxYvZQnZH84endE2gtlNT6i6nglkFNAXM4q2KxSFy/Gj6Kma1oPaoxGx25zLpZ
Mv3gEqpXoFO+cb917kmtgZ7EpUanRz905Y6b5Kk4qUjI7kyqtEI66qvTjKWCDOOs2qfEi/GB2RvR
hg17OZ9eECfYObpb6zGm3Y8+oaxZU3PgtUbJBCMklgTFz6oni9muIL4FIcs2bMTGV8pqYeYeJ/m5
U5AWlazOqg4Hv/zwiP+9bgGEZKLI7NiQv56GrCcHtEeWDrpD8pspQkf9xz4/sAw58VwoxPg93RzS
0d9fsUwMoOXhEkqz4sxGofvRobKeTKg1Ujc6wB6CAGDVyr0Vt79bRydwTqO9F0tHI2K6OX3r/hQD
uND15+1WkabO1KIM6QAHRIzxogAM3kR+G4hk39mM96pR0oc5JzCMpbpOthTvpXc3fsc6XpcdUsi+
BrdQvE6g+hQB20c34YWRnnX7igI72LkoNBuoG6LxtCzeC5GqOuuFA7Vdz1rdZnhMmAwvuF84WEMl
PopODPDyg3ICpxtY6xk+ZzrN5p7pm5ybt+88GBNa57hXpTT4lCUp6tHRNz+1qMkotF7HRfcqL63z
NQmQ1VJXRISu/RC6BrveAkGJv+oMPZtsowMbvVoXwBbWDDkyn55q1pm/4csY3jdw8jnUIsTQQVw/
2TOX3JuUNTDccvlrnclNdvv2psaZBn2YmMUh5iOW9cIju85iab//LvnQckpwNolyyJh0w6Z2BGtu
+PIzCufv5chH/6JYrNoUm9BCQ9V3n5hwsebAiSOg6hilPVchALdT120tOMhVwCUEwLOTacj72/nr
+DSmRHBWS2huUJtidUuVqkCznkYYzcVzQb5I2l17WKXw6RbfH89beloZ0FOhJ4IcfHyHM21GII6x
nDDof9nUsqAjoDnLcPBplG4EjiE3mDyBiv7WBmJZ2NiYte1ZrfQ39M1u0AbOUgbIiNiKS6Wm234x
mUHk4BHVQUBhfGkmbYg0yH7tlYoOm4AEbMLHMoq89Z6GtQaMkbsGG4zRxX5PHPPT6xk+GlMIoH4q
o6nAJ2AJ1mYmWLuRvtF5wMOfDWapxow5gcm8LSjycJ112IKwG6ymh7e9A2KWknDEzHCGr6uGvN4X
7uspe7OwLH8FO6XomSOHiSoJER7zW8X3bVwI2aGgIIqwCb9up42OpYQs/z3ed9YISEsdLfpNuro7
uQpZndBxtbI5B45k6+9U+9IsDDptjWqYA/cLrcMVlWePtQQW/Wvlg53HlQxnNrcwnUEF3HuxocyN
wWC7i9msT7975MMzeSqKVAoS4rxEkpjjOmnSyJuKWJfL28sAG2FDdRg4Me6GqgKsmqb+cEMh0WjO
3Y83VgG6sDZBuj4hrOjw5AQVm2eJ3bU6d0ce4zoUyBiIwn9Vb9TqSG+BjcWM9BBpZjztfDD83tur
dBCbIs1ZlbyOTJQTbbqJKTmQ7rGPg7XACNzBfSYG0srag2udP9FW8PDHqj3hqaUt0PaTurf6iMBD
IReNEGJROB8m+J7QU3whfA4knVb9vouehxPo99KQzUDvIn45GsxyJgav2kSRq50OktHGa2HuzTwR
RguB1en/ZOpP6JE0JLSq5TJwjqlb42PAqGT0P+pElUQtpQRLkFoIsHKa0iozHiwkLGQk8zWFvVL0
C292Suq+n7CDYztCaXKdVvXb3S80i/0OAY/ke+PsrM8GCo0xLu7+qTYNiMdcYb/zwIqowob7wNUP
DqBbcYbqBl7kRhezKwTcFS9uppbvXirziZn+v510apcR2vfq7SqLf1B9zb4/9dbDbZJaofAp++Kb
ud82aQoXvrqOud/nzG55mkb/v4AnVLQxIo1SQGa7lzXrlineGMDv7llexZLS2p85zlUw7y+wVZ8s
h0JvHfIkUaYQCihni5Acd0KRzmGjM62ETJn1vloN5fb+uvyySNdcPJDDFT4GaoQUVk1+wiWocs3o
zMN7omjKAJ4bRKkRjRXm8I2gX6RVjIxEZdeDVbxpi2ldzM/QB1c3s1NDDvW4mjdYfbe7ZSt9WkcY
ftOCmgH67EhCuzCzq4TTjGqiDvu2xVNwQyjvrSeVav0Bha47YqEDzYAY8Pm9FHgu8RjD6gvh37ip
63LaiNhAiR9ZCnQ85tzeZAlqvtOjcwKjSqJjdzu5/pr1iScBm/nsyu1WyPILhKrXbE9LV55nmNMC
cBSrkxgaVyaVxt7Ckp0OgN/0JQodxRkurzJVd35m66n67DrGKZIZM4Q90/9Ypn7eJo0AbLR1pRYx
bvJSKmGvePfy2+1N1jPFvKmL4zWgXfwi0Yzc1eOUpmHi9B7kLDL39gkRltlqpgW8nE2hHpxG80QY
kh3e0X63P0m30TMHIuwu6Ze7rLz27SvaJiIqxcMZw26JoPHhaKlciUckXH9G8mlXdUXOl7eu8rSe
9NkN8l1HadxZexbeoP614yFWHkerlD7nNto3se4xsyBc+yqrw8ZCPvN6XiAIg2gSM405iHEfqcdu
8A9ri5PWpqMend6ZX3Lx6QRmohyTIjpfT3lgsThdbUp3/toRCDNKfo1pEY6MlM7raxr4x7cILH5J
q2fHJD7rtfjleF+53tH1NeLUOq9e0wzZh/d47KrfZPbOQuXt5Sgx+JmIL9u86H0rHp/Q4pt2BKGU
/8lw+9wghQiadIqUJ7UdzooK+3ZNMgPgJQvNQS3xwpBo2EPrB5dOlBi09U1+5+y3QgZ9LXp9LMpH
POWyhDNjLCA5/3sy8eA4ujco3uAW0E0u3lcm/zom77U5fUgQRt7tCu/4/nQHJ8T+blcKlS7pnbJ9
g+cj6c1jLFWGduQcPdsFufSA7wFcS+q7yoT9xfGfxKyC44cVH07jjWqgD/RKntqsc+sPuw8nGwYl
XWitCjwj7qGmyIir0tmlxSXBNUJVuHou/k7jGi4KQZz06HNx7YRaOIibrvjGS3xWRI8+XPCvv6xt
DGflq5IzB6ZdJ9eHksZtpub2IBRCU7S9PsM0XMUdJUfHZmvzvn8xHUwPBXyGZwwezA4z2ay9MbIM
8e86CE5jp0Ozh+tGWH4hj1EGzjhcXOgC7vpU5JdTltOMcLZYwKCGlcOKuVwVJoS5dYY0qumBW8t5
4hyL47XYe4tZ3DNIS4zLSUxpSu1NZg0ZZUFKoI7QdT//Dee7NLKMcZYmLImTTA9TwF1TpdxqzVrA
LiKYMEzMCa6gR90/zsXA3Bpic2gTf7bURxyaxA4sQbtXYktyZU4M9glrBAqQxRYQqAiTxt0V5F5v
lS0hpv+4d5MlA1LX1u0blXbAYSDWHAzB7FHK4nHU1lnhTpvB/iy6Pjh7NA6KJVmLihjij5sJrujS
jpUC/ZGR6VLex2jo34lViaOOp0XDV8snd1YktiZGd0uAdPLr/bNAkpTleo9fNKdwEdZEODP0hMyI
gPQ2pJ/jZghRQ//ah0wZscS6NAcS7tGbTerqaB8gL5TiB7lKcBc6jNFMh1pqpO8LqYz2DCgPQlE1
axlZe2Z5l3VZR8HjD0AIDTBO297sFrcECHZAKrFEz4HSl/TZWs/cts89DcA99C+MJK1yJQpGtyc9
zT043LDsntGCm2kiZwE/zpPhWSk69yQscYNkmPEdb95z4eX562f2yff3OqzaDamZzoO4fpx2iuDR
dMu0Fnvnqmr196h/rhgGnQ8K3f8HG2QHRt8gDky0q8UMvhS2RAK+4LM5Rw4itX5cnw+qCvXzhnvm
bSJoWzGj2Dv2f+D84eyow1POhScEBDFrHuV4N5HaAtc8pddyBGdmf9nEylkiDQSqMysd5MJMrBDd
Ew61q/KPyzsNyy28imZkoTpNA03tgvgVNqnRpnEIIfQTfHqnjZ6QJEXWeVo/IKY9x1na+Y/SUl58
s2D8110LM/7yAC/HCjtlQ1qe3o4aCXuru5/qZ4KMzA9SuEIO3F1KCXg+yxMAX22rhT7dyHAsGHUs
cUzRwISbNLR9BkgX7onYiE7vcn+GENoPtCOJKev3pWOoWd6VXnGxXz/l9ZTeu0LtI+vaU3sDsgwn
0k9vC9G/nbTnJ+Fu6GIwgeVAgfXMgViadMcD0LKzQPqqhfg0nmBxgEtVTZYN2Mtj91Bjp8Vg7QjT
G1WN906LaqfOoMD4id6RvK4qV0AmkuY1WayUByA3PubbDtt8diREvk1ofOabTKSOX6KYmJZ/AMfj
+DDrSs9KjVkI9ktakwZp1uuvH6A0BS9Eu3378iWayTcUSvDdzdIpTYMEv9fVWxnl/lMNBgI3Nyga
bE3CUz3f0HBh460U1A4DjidfgRrBJssNkSh3uS5eLJY+bHQBqiTCk/YXtzh2QcBfEDJcUycosB//
oudVxigIOzS4HHR5/MWpCTgMhtgdKNrNjt+jV1GHu6uYFGcsb3MxpWQXKvINUVTNPEZIW55tJ7Jk
HKFD5H3fjL3g0uIG9tzOOgA4/GGtz0lkekzVpUAuGo+pYobWoU9EYKk9yMA4mHxpQ3qpsKTOwEdn
Blkfk9dlJFhC6e/BZMQByRm2FFdw2oZ4q0zYT6TwnIkHk6fEYR7aHnKxffZzS+wpt9wkVdLMxT77
Z2V3B5VYBRVlTqT37Hb5nMF1ziyUuvJU2kqllTpCGhFt5Mj67m/G5htLv1Rh9LtO6jPdfx9qkDt/
smQFz2weUi32mB9U/c1zQ23c5gBpdVpt7nVpwLEqUGwfxdxwKEaQEMKPHLJql2ATZ4vXFeKaNnpk
THC3VqonpF19PcPw16iLfeeu5p9CQ5Hau3ip4WCa8JoaE66LvNtMm1oWBzJBVY+obJAVlrukIWxQ
XihvoBPSbmbkOU9pmf5wlpubbwtm/5uAeVk0MTJZaxXroEtp0HP6YY4rq2tooflZAIMS80ghfsQh
VbcYuVh0swgM3sOzeqPmZHghinR8Irnrhv3PNp6q/dW/9NKtQLcgaBh2dfmd+b9fgzU5jRtRxS//
mU2yJKD2HycLZEUDoDAoE0g9nr+THa7uWNpaROO0iORW3Q+/yZzrnDhBWXy/+a5Qh0jRTFKkJPVW
TZuUxmY2uU3TCpCkSBJ9SCtVDHL9W+vT4+AJc6/yhevZ45V7y8S3JWcWQu7m+yguZWevziyKbA2o
4157evFMI7ufK9laBvDsgczrOxDzMIiJ0cV6dMZZ/c5lKK3oh8bfYC5I0GDODyW6xb9quxIGFyXp
3PF7id3O4KchmaUNBJdfP2ssxaBNkw0sMlVLLUdN9ZF4QCgYVsHLxPcurCd5BuZQizWMuc1VsqWq
f2TvMKkwbOFSF3fGsH428izY3hDMcFVZQieLyPyi1QP3LdNgnVgDKtGGhpQ9UUUAEI1fypqdHi6W
Lnv+8/Xb1Mid/MA7uEnF8KdVhVze6GrmbS2kboWVs+phcE18/q7ZAqpIeKByiVuwxsg+Er+RgreD
8sgu8CGVNPJHujN+uGoLq2zbS5QDnEiokoS46xF+bqCvRzSadxaR6XrFi+KxJDaBrtA/6+uhRYVn
vO03aT5YxdKNdkagpNX6lVTMuIGxr/3yCpaip3BRzxUwbv3CRGO0MhheL7GwE1e894r6GvUiJ00H
+qnPQCXH84t/svzA4GjqHJ+bEOXs8alggtRHTUeF0UKm3rhddds0oz/qaUy6iRDJfa7hyTg5kXTf
fsLTdQBGwryIFRD6ei1bPAd9GsCZpIJeEXNFSbi+fAKPxfi9MxvcwW3qr6mJMJLyYnMU5BLf62GT
5YMq6apuCDMFh6B6TlJlBMPqa5ftfvCGtp7bGE7AIYHA8QNyFaOv3+8ENAum6aD+AEjRTgjRcK4S
tgs7rkxxxHo/g6xBo8dreFGzcc3q6l6XcDmNTaMP6lcjUdfUnNAL/ZJCO/pPtqMkaqo8t89kKcSh
gUfT45ZIy0eeHhENjQehDA13LKpMVgoIenhNNKpLRmm54pullt0By3h5Opb7wsBjiT82TX8fRDnU
eeuU3hh33ZD7dcUap+3gNFqWxIkvdpbk7DK4w0EY1JXcHXPTSiYdSONmBZkj5PyR0GwThnr2V5T9
ZroBARUoDTy2fLXc+IKatCQWpE20Zb+Xzzhp8Dud/u+xhyHWlh36hz3+Cpv6U9iml7ubFEnNBxsn
KVPO1k+xlpg54wILB8B4tGHUd1NmJt1MkoVx974YJhK2YY+9wp/8aina4Neask8q6KTxl2gLofS+
3O85US5MdxvJ4KUx4YkBMsOWQj6q2GXk3v2MJdrD1TcI8uWI1qMQkzoTMbaGIe9WHj0xOIVOsGZR
kaKim1d76reHLOvR8f4XcZgR0VfPYyBOxDZwYklZ7zc/y3uuPJaLEtXxkSLcOez2NR/meyj+EGpF
qKJQ313EbGc9mCOpu7OFBpCDcDw44ehLhuiq1vT+I2aLiy91nS+h1ik+knpxq9kRqmX2cWoAXBgV
WVQEj9V9LSR2/HHdvLMpReqI/PHROnl8f7QVHAFI2V0cwbaVRkWmpZ40H6kSfXP7fgeDO+tBxQkI
npmUUMLPSZHXqQK0gA/wE5HHv3YMrn8KEHEzXIvlzUqPHY9T8cYgd4wezkoJPVCLQ9nVP/RfgYmq
6qP+/06CcJYf9gdsi61YEXgaZN8GjgXWstowwrKRrX97xg9dlmCZCQtW29Bw3e1me8fZ8QSy0YOY
gMOlp2n+0HXDHItDvQyulBwktNJfcAhyAa5ZVHkZKKLz/Eun0gip88BgT0iVXJ9A1Zp14gSf9zRV
V8EpCAO52PdC/TVjeokv6jhyw1s9dW97x8GxW6S2tUuWSwBZ/rdIr2CYB54nszTCitFPRSTu7BWl
7+9gB5TGEiac7ALslCFFv9jEQltG+4tH9Sk/7/xCXyeelP2SOlKHIwWo++ovRLpPo4+ztxTjJ9hT
Xik0DTZmI4y+qHSED+GTk2f9VZpBSqSn+F1mkDgVOUL3H9ZFDka7nJ/nTC/vqlvsoET5mfSu2o76
MckCsFyVjpPO1ZOj9O8zs48M4lrQinl1JQJNo8v2kVGl6MuVKOoNPSt5Dy5GDXUcZmyF7A4VfzDe
jgwIrDuo19gim3YYmZncf62oP+1lFJC4VYR+pkUasIQpcDxtBjOziHWLUj+dCn2fx/orjSwqzi/I
Wb1mOWpNY+YOlD4/15h8YZoW91vBmJ9bhjV1KMvVDm2mp0OdcK/IuVCpLXJrAS/QriK9HehlQujK
g16LvybqMkoxXbi1XQZQ54XQb8RqT0KOJ8G3r9jw7CkD7+btB4e8AbVNf+YCTZriRnHvCtshNeEl
NYyZ1BD1GvPD+XRtP2SVl8sIYjSaRi/tJGvSYm0b8qPgkLEVGvQYTxaz5x+xvSPOm0JkVDCATosp
NhyEcmTic/W7sfPO+SphFJicZNxiTwkHgqvX0YDe+rZuaCy4ogJL/jibtZN7kOuGl0CTaiLzF0V/
GQulMx0d+V82+g22cmosijeEwXPdpZSvDMG+7FJcp9SVCD4z46/KrtYW8BOKAyRqkotHNs4qBPbN
ERqTIs4tcfOqAVh3arka5/aVtbg3xffmJNYTQguaIQqbfeyY2f5pSmA69H0Mkfu8xjWnyENW7Ny6
ZZA4Yzx/et0ToCYPJRxahUkJUsr64LR8sfijLvkPeM8ERJIwJTHKcPcDeO0RSartlPIVfqOHFoqW
jBLW/kXHFKQZBYm7z+6lheeGskjvt9ugO5FkWbiLe/VFSlt0kMioEq7AzzOYiP6e+2o2SpJdnW0n
Nl0r/+ulVcVB6Qlh/v8K+xF2K0WVNgOvk7whxGChT40MHYmRD91wsWleKAXWHr+yMj+9dXHICBCf
nFLxISu4Xo1rmJ8pbDiuxjKWqQjr7yLG2JekVUj1ymT4tuTpDYpc8rRWe2AnMkYF+faDhRaEzwXf
u8m/LkYUDy+p3BrdFlaonZp7uBPzGkfhWXmH+p8SlT2l/4IuSMdp12PldsCzje6KS+hwwzRvzoRn
f+ZoORpo6pvtUUo43gw2akQ0wG3EFvU7IKZnRx9Gb/9cgeNPp7f5/3GLwBAPoJbsiglmbo11oyNA
L9e0oeTTXjZKZkLsLu/pbi8A1KNdKskEutE/MzdYgfqU0BRPCa7jKLG47c2adWq8T5TsV4Olc4KG
SGPnNjXV5ZNFKXwxBQ4cWjO26BI1YUlubbzCX9iXrt/m8JBPwBkG0Q3WtjjfbonUp/jC/QkU/JPF
g4J1pSU/a1HJY7fC9/ffFrFSZNhdejw0BnHurdRIs7Jm2LJVslZW3fF1Ux4R3JCMyvxD8jXND49E
h2py0QvisCSE/52D5Z7om0KsuoVSBiHSzb9uYTZHbGyOVjA3wEcKeEdtiV1p/Sz2ZKwWCWeqWbEB
V7siZqdkr5tzaJcWYv1DW92k9FvCyGF/5PGdFMH+hZV632O+CpqImVwX5dADmG73nvz1gs2oReeH
D6JT6PvTLckP8jLS3xbYsF9zDNK+yvwnhSyLSGWZKgiTtApTGbQPgfrv5rZ8+0Fm9VWU4tONxCtG
FHdUVSepkYHeqZ510NbbUGHlg/rqDtfIT2+ISgjSq/h0FnIuvo1n5GNfKN/jByHjzP8bbTSyFVw1
vgcdgBEH4XK30hhSEG3cYN2xBpi62V9gnZ2DAlz1zideZzA9j2zO6jqwMz1jCOGYTmzWoV6N/q9A
Awe0L82sgiOgTaSc8GmzlY/s1drJdJsoPwL15Jrn58LOHTQcO62mgUHczeO29E4a3wqqxhr/CYZA
ezhPIy7eFVBoy3zBf80gKl8l7P60IppxR+a7g6a9o66ldeOhmVp32Ol6Xq+j4/VBEKWVy3lqZDZJ
aIajWM1cNsii2PHrSe9+4Z7qc2Im/HgSWvOxMgJJuP/GcKHMXCeuQ9WSbt/74m1EY/3Z+k77ailB
Cbwu4vOGJQHyYGkS1DZ9KZJfTZgJ3uspW7snILYjhqIuyelPqQ73GsAkP5ZEYofKO5hCpp9puJhE
5FYjveYnwvDqXdChTCAJddvPqemVJ1bjjxsjxdvsqF/9RwVQbFHLfsrx9nxayfzqtqht4FNRB8nO
bwFVeIUgcMqDgs4CKm9MBeCF55yE+/GnCTEL9hXviNOFDxU2f5R78SYzwKo98g0Uop2HGBvXQw7s
BOBsfssPIcGDc+3NuI9gLtC1zUw0c15lyU8CL9E273enzEwaHOVzdvflF18LiwEwwHsxabQCuj1U
X4G8iCv7vSeXGllE6+Go+wJUCYiuU+Wxc4/WGqCm2QCKTqVh0y5LIJVcWgwskZ6e7xEf40t17ioc
zHND8mkzzSU2xNGcvDdG3Qh/cbrEBQcPLKAcTxFMKwG4K91Ih7BmvjP6V8ns9d4GCIiGziy/0W78
NWQTP0PPVes04b+TBnlgcrAD3SsBS6yhQwQJBRd5qE5CKuUSGPcSUFIGv6cFYwhBfsDrUBP0urjb
kmfz3r0EfzC4gBT1xP4GVkVNdDE/mSn4L1qSjzrcnNA6hPKFz6IiJlTFufz7/7uO1cYXxvyv+pl1
OeEGG5a7MKLn1ZKFWFMQE+J5+9ZUx0XLJak9sWb3gYxGMhBCeVo76Ik8pDiwAIoWGRLLscPkXKuq
dmVbw64Er94MgEaIoV3+gKjb2chUkDlw3HXYWcHDtOODK7lQ/Y1qMXdECx0MQBpl6GwHFriDxRd9
9i+hhjZ8jbSwUwIxXlzAGkxINuz3qHRJTIgJw8pI4TqVtMAg8jZCyfagEq5PLFjl/tUmXnXPbmpy
hpPu3Xwx8udTMCnQKs5HPYFC/dBfG0YBalfa1I/lOJz0DRMQyX6L/wpsWfrtQr8zhc6QDsx6FFMO
OxRDVMG00+RtQ8R57uKe48ex29p7RggVBs/19CIwwaM6RRIZ0acCNU+fYbVOZeh0E2rxeNf5gK+O
v8Li/38Pvbf7R/orCqMaZznT4fgVBlyJHd2Dd+qY1+HxS7oyVpElIa/6K98ICpKQfiZa9AiqM9YI
akOeHUmf1Y6XGCk5zZE0HpCDMlnWr+5ksYgYSeMCoCOM+XBsNQ96ZNR1PJ8Q0g+SB69chsUV8XLR
NXS7kcVuziQArdMaapGIHPJVSpDkSkXnhjAENlz4aP0IreN3kuCJqNRuPUqYG3rH+up7xdtjAJcY
hdEee1ONqisSJBVIoTiIInNrtOkYIgdiSqmQnUHNF0l/xnUyRkFPwqWU6QN9Q5xcjmCdUeKwDAnU
qh/vTB8BlREG0AzEWlZKizCIEshv96nNI/7UhHaR2u+aVdFRIguuhtBF/Pmb8H/FRTkr4FrH/C+p
Jss3NsbnVyZ5+PMUzlkgR+Alc0JOiRh2pcukpAfhjdMn8oBf0/2RfFvdO/69BzXbkBkOYQjEobys
E6vLlonM4ix7MJCDVMj98ZwNCiMvEQjj5jJi8RtfOpfQVcIH6naiHoM0ZgJkw9hV9698IRsgkgRu
uTq+ewOQ05u8/xoNPpRtF85H390+FYDaieU1wIXM74oABqF7082+QlWSS4QlB5w2tpvM8sQZATCj
kBq6yrYATF0skINFfryYxQhK2/tUvQUTd08pb1oIQjA6oy6swOiw9j+Dbz7KVzUGlSnmKnNFeOSk
E0OkH+ft0E5Jgaeut+gFJTeIb6HMdiV50sb6ReGRJelkyHKXpf9sVfQpr3hruZEXnI4pv4Ah0oJw
tGTgGIT2AFus7m+XBHp8+UiKaL984pVUHbqbZngolwEJvGrtHmhMvt1G5fFRncSN4YoJzdYTBqZT
G6ZRgJI93yyloQ9JjJ4aNQCeT1bN/tgulQeAgQaU90V9QAS1hjDLFNbIm2l7pleKXrDm1K40Bhkj
F49pzWq1xGsfLzZS7yBL9UbdwhPgI7LsTV1OU65bUlUod+ofAp2CHJCil4X/dMP9/bE2i+Psnj2q
lVxFTbvcTBT6ds6oiWzktKsEQ2tzVOZsxLE05WB1W7BX7fPlu6zA/ISW+GNHikLYxHOsHJydFFtS
6rg7KP/jjoGKShOUC1Yjr8H6idSACewhclYMZEeHR79Qw/j/Le6A2WF6YsA5NIySI3TPBJJAIaI8
jSFZi5O7uRQeEoBs0x0Z4Y+oEKNesNNcZBSo1/tl1b2d2A82alTrnlw5nH3aJIuqC+sj7j3L+uyu
U7DBFfapQngELZRUMRp6CqMRwTe+V+aBn3I08Vb0KQtD9WlL7MDJl8El7E8G0EEM1pBfcetPJGa0
OQQsBU7CtEm18x8SI966VCoy+bFUS9PetWRDRYCzrM8waJLtlTeEfwau+vq4zwmZ2YKigP1kpCLx
2yfpSik591P3z73c2j93gADjbMSsGCxxe8ZpYPI0rD+kvx7dFh2Ft4lmTvkQzWiCpRlvkGwR3a3E
Cxo45peBRz2zB6aNiPAmRCN7rW9X4VHvzMuP40hhhrfBS448Aih+h2/ysqJNICt1bsZMOK13BovY
YFZO3yb2jxOjgP6M/h0PLnXdiO+qzyfjRDWAu2do5tf86B+LXP/mdemrmNanj557SL+XTG+e5apd
uS3DHoXeMMtW3GExhxQ2Zt8tVv/rlhhDcEfqJLku+fMEXCXzjvOOsyrs2rK7uOyNLaji3aOmUJgK
/KKWmtOHSIQ+jEpu2qk5B2MwCuV1JODK5ZTdouRKrz5dF/pxOIr+2xoQMgFUmlEHE+98nxdOflfH
qtdGG41hCNHGcEXNdgm853Sx7b9Rdc8Mb6lXItTAIlarEUMSf1DbV7HuMyU45oeVCX8tuqh1Dl0J
+TPM/PLlKYOURBYUMIALNzfNHyYvMTrsJPKHCJgZOeBXeorvpFEx5gMeadMmJUw3IUy2q3ifgKNE
ZiwtE2K2SvB8s4JbHdqyqqfW4KyZHNAC+Pg6TTHbrPCZxfSS8dEpGte8mnHa7JDsyGWcPgv2mN4y
73OI1dNGfq0zosWQtCcMmM1Zl6rSq6mxSbbt4EIj+EC6WTa/U/3n/0AfGle/nEx9/5GcqYPsO2Ni
xE2N3YVeMsmRcM5Mlt11CH7cRLI6d3Ne4fXAoHijyzyp7IqiNdJ8TgjzrwxdxkXtaDvB7S7XyxL6
ybtk3eKIQ8CR7B55k9C+4A1KFGrkBiHrF4LWr3k7b7gFUJOIW7NGAx6SaMilJK5lPpj6eRvG7DUL
uQ3vS4pGp5CwcK8piSqEE1nswAL+IqoADGWy+68PU37NuzANpfox3/R/QeLtyJHtX6umcEVIEpqa
LFR6+uB3ArvAr/r/MeKVWczowBblWwXYICkvjlyWSN1hR5SUySgb2sFwuXPo7hnrc/iWC08sUx9T
xTUt165WoUGPJ9Tbxwtq4OewQ0eYueFhjy6jL2BAQNpxNTmy3fAS8A3MlwRxGKjsMtDPziER6muJ
oCRpcyXhxtP/m94y09DBVMbHz2fc2IYzyOwRCM+3LNOn+qbsEeEYyI4T3fMqMDi82sYYYKudA9+E
qrq5zQX1hNwPeICZeLBpyfQAniiNEal1K/wRZvpP2M0X9CC6PEw1C0iBYNrQyMCIspUu6rIi4v9o
zw+6OWxCD0P0Xdot3IupTFT6VHIxY+KvXiIyzYh04CkSJ5t4o3C8QWCZPlvepi30xmE4f4x3P+gW
NihyLOhPku8o73J7Vhx1wLhXP3zbYhJnUNBa0QIuKMoLfGHngPCqj5JsEgSwLXkUv8dFXJy2apm4
rnFyN/1m+oT+K4mox1QYLSnqDuBolOyyc5Y0Ia5Tvd5pFwqt2TJ9mhoHB3+39Qb0d4jjpr0Z6m3P
hJv8Wjv/xplhjVATsRPO+N/H0SzI7Pd/gcENDCOJ7YIkPDx9cPwUIrOFYKPvkqdnJD8PI34rHKB1
/AgKywHPWPeqeLcdD76fyQy2rPMUGTapnW94ypfLLvfzlzj/6quwMhguJJy8Kn5kh5Ecu7XfrfZj
abrKnVpL08oAxVl68dO66ZoF6NBAc2BiWWqkqhqz7palWCL3S5iaqfEvr0BZuWgPYomiXWZItKHQ
ARgl4UdwLYLkWWLCJFJflmsMY0/UbBRuasVJdPr0V6GigLnOiofeBuPocJvqVAhLSlzQ3padeeoE
i3VQ+pJV6Z7hkKqHLd6FSAYH/wX5hZDIynk5kw9ZrMuRCAFKFSv5aK6UMBAGXyl2KvuaF6fR6Ezq
v5+ebg/fJp8HkuvfGBdWp3c4O9ttJ8Ud+Bk6LqhqRnzW1msZfgyrgUCQafzNK+MYhXQvhO9GfC5P
UnjZGp5LZHl4N89vSpnqqOq8l1Rzk523HD4FZngGKKlbroHzuaf8JSVOXHLRVUXnTj0ZOjgeDguK
HgCWB8A/oVyFopfxPkcsivj1QZPs6k6UV27Ut9Z+phs6xrjxep+euM/E8TMdaJYS7AoZ0TsIdNub
pPWWX7CcP5cElZhjtvlO0Uyy2bYMxqmEyaPl11a8cihgBhnSaOboX6AViwAPOPjW0RXpkoMGxrG3
naNR3hEwr0w/IuiV0yjqq1rOm+nQ/utQ+X7oeQou1eAu2XfEZBB+0NI01/dCUkAO/ZxmaEcqJL+c
RsdjrlAE2QlbvW/OJVmq58mtwFzJmEHheNJBaAfwjXCwe7bezQ3B9kuLbRpskU5ZbqzpRA9GDw5Y
ijS+Ie9naWOXliI4bR4KKfUE+V3+iHqmqNf2qsWN1wQz2FKBwKWvK39e7ZRY6SmdC5cN9940eRkc
B3SnLeRZl2C3UDA/5kRr3enUARrx9SK/9J6Z4K3u9UY92+xW2lN23YfkoIe6d71eQ5qQdnRGK1Ek
OsILld8NhwNdp6A2qZ5wue3aAhmX1k0jQbRT9/hljXw4rfI+hh2AGJdwYw8YldOE8bfSwkbxqb1j
+IZlEKYp6tmZsvhSMMtEwxTNfW9vYQ+Pii6+n+3IevClnaJSJiVLp8f1Ue4TrhMiLLDjKQZDTCZH
JLnCza6PoPgSdatLffCsMbaRcla/StijC8+eehq/BmyB5SrXyEQva3n0s7BywGOiABTwWjj0E9UR
KhpmgwyP363oAHpQluCPx9QtMCqmRhBM7bebA5EyKMt5q/2s/QWlEq5RDiNyKWn25yczxO0Z55fd
LAm/gGIJkS55gxO+36lmNER+kBr/9X5Ghxr/GmAUCopAW3GZN1unS4Tmv57L3lOWiXoWAk5uCjeS
b6JWFwRL3RrQqbFJ7zH1ZUMz+9U8eG6t/XTBl1Q6nxP160gX7vM6Tj1fAjC9Sgs1c0TkHK5Bvz3z
IG9L9GDp3uELINLwRTw9tuaArNCz4ujNh3JPM3rpTSP7b3e+EqsOXv1O/h7NMNWR1de3TgTe/tnm
T4ykPtBVJ6laxqyzaQWiwdO8ML2d4UC7Kz/xvcfQhldDZ8pmkCuhlQ8QTSKYrVYM+rXuHGfnLT4f
YKzx4YjOSQvEdLaNG7z2DNt8/wif9Dev5uyw8Rx1D2TR8nZyMJ/ZO68LvfUgugocZ7ihKN5/zctQ
tfLj48IVCiaqh95awQSoisiW0Jd1GvVwda4kTJ3JIbn1FaDxkH6vnvqbfh5ChDRLID89TOPvjQsg
H3fZ9i5hfykQOduaDb6AoCeZS7D4vWcLhiMeiyT8aphXuVOAhuF1VwKVf1H2FkrAxhamnBwhtLht
RwUEl9jLpaRt3ns51g6OrwH9gvKwqa3wx3HTRU2f4tSl/wkYyjtbfX+M8Gtayyav+j58CwRXmht3
e+CgoLVp86vNslqGGCHPpZE2Kwz4ctnehe4BCdO9b4yu6f7VwwaJCrQAVZi/elu+VLb9vLJko28N
Nhp3+LVJBoZOoUoKecrQNWFcJ2xfshVhVhK14xMd36WDYwseoWHjrTigZcqQn3bBffW3HBFHj3G9
SMBOax36jC3TwOFRQ9rbZq4DkNEAKOape5ysJU10E8e7/7WTBk9vBiV/r3YpXGY8+E+em9l/EJHX
vip9fy1Grvu5at5+zwfvvgUEBemg1/iqhxggyT0zup+dRVMp5oKq8Yrvy3KFNxNzujVlHjo/ym3e
HZV7o7qd4JcCFi36gmXxzERf23J+xYRqabq6uDQUWvd0qqjWUofW/j7G5j+2zqv+uDO8BI+5G7tj
65ELlGzEzQHd43mNZOL14dyJLee2ClOEHG126vNz1TEW7yTe6lt1xfiHV33zJs/DbgJHJ9rjkLux
Zcg2wnMvSditcxGmGNKqHfGP/gAfmh6CplVCfeMfME5+wqpBEW+PldwjONtEqiyl2n2L+6OvGJJu
/50chbSKFRTJ0RbJeoZW4AZOPeM1FfJnigvSmpjOokwd0oVLsmj4fAfsH3cHomcMVsWESrNoqej4
0ngcJg3kTi99pBE3mmc4nyo3rIE++d6oWZ7v+MeehjjyszpLBkGBOSpZ8qaCrk92tPg8rXvki/+u
iTOmBEEIT6+8HUXhS24aBK+4khqjD8rveCnFIsomSAz3NVmQZvCh/74vnYZaKUj2GFUpjYctbcq5
51lyaYmDmYLjJEzjPaWTZZBSU6WE+pMUIEAZ1KXf6uRqfnayB0zCurJZCv8t1SZjVnDWyJXiyDm+
aHbLClWfzXoSSVxdlEsZlMserMoSVFjRHTTbg1Uv5L7Ae13MB0u8T16aO4aBHwtXHlKFh4Ko60XT
KqpUilnOtI8PwKlRJlWMDeBbJdQRbKN72Z3Y9izkzDQlAkOSPudoIMwutToHbAFD3Pg7oDW1n7uo
e7SYL7nF59ESsov7toLhhDevjvNHhDcTTD6hgcjV5j9+VaZnp+ru9HTGTN+Ni3S+u7/9HyXCGA2l
BhBCSJPaCDAxhwOSPOICxtnCD+Vm7CUlmXNcPxTxVqeT66WdJp6u1J6FJteZgucJslP5OL0oCdA8
SLPdVT8z/jEzCZKEw6l1dRqX0ejtMBFKwcZS/o8IVIZ44B/HvvcoVa9tNcEI18Ht+NgAgZQcPHWP
TgzWPJRwqT2G4OdCl4ZBztWf+ANi+t+FXvzAUVx9TP11QFuYlN+QRRa5n/8vvlvxmumZa+wAdR4j
jwMWJ15I+Pkl/xK5hQuEPF9+2LTJCL1+v6lvsqqaXLHXUw6VWrDmNP/Sh5WwHBID/uxXHZDyz4Mo
BC7aGGfgaA+bPBl8MS+N68jWHVO110EUgZgvmuRgRK2tTrAaIgrzB1P7enH2QBiaCzKSWELOADoW
lYG4UrxwDwgxy5lIl02cI6ZsULSwIEGBJHmLiiX84Tossb5dxzdoKt+EdKyZjGQ1hO0NvZV8Eopu
5jqmIYFdH4RV6HDq5Oz8IrIzQbD2EQobpIg9Zpf9AulfAng6ME+cNhV+fBbJJ01gCJzNl/EbeAvi
te1g9/PD84y5nEJoSTQwfBQgiD/F0NuZwC27Qbeh8DYsxtuHqYj6rL6/Hb7+cGUKPP+pkuhfgOkj
15hBPdOA5QnAiQwRrJWlpxzqUuU1OLk6f8P74nHpXNdIi3RwpwOe3pvzjdni5yK9KhEjvgoVo4hQ
l3aaW81en+TbVzr31jWvJZmqEuG/IUE/wMWyNSGWbce5NX3bAoDAl8kYPaibxn7Vc9W8CpLhLQLO
RPPPLNpd+rdzvkD6NxpjkcwdZAWsAyDJSvZhMM0VXc59P1tAYDwWBv5jeDk2PlV1zRh0kF5Th/lB
3cIeIGmGdit/6WMlyx9EpZLcyoM1jw4GdH1Z27c4WRf74bq/6eZhN+MDQ3rTqmSq+fJOZa/39oC2
QpQTpYm9Gd/l6I02z+IesmvOuglEU/2CwKlJoYdIxCOZMuBnQqwj8SrVnjwtykC5wRjFukjT7SxY
A/Sv6N672gD3E0c621ltbqpz7RGUo9Oam2reUroAoPBMg9k1ZH0cAA0gtnGPfMiBtzknjlqvYjbC
wWUErrovma0SYNJuYcyNd2mW1BE9efvKZwoehfPkBPQKffLpTO7TRlh0V6y8rwEBkcX03+mxiCBa
3B4m3hG0+66L6+0qEGYMuezGdm5cKpMgqPYR5dcxzk5H+RtMToo+RRT88yutS1cDUDhKes2IPLMw
LPk0bepAM3XmFMq+nVW7YgeC4AHGzqRdCcSc1jaaTNV7IAnD93k/ztSpfxvoFTnix1UhezpvFtp7
fDNtlNcowSpsAtENt4EdnC02oICWWs5sdX+riWnKoEg0OSh+3KkshH/HDYr2/C1oOONpCgTM3pim
CR0/N+xrtcb/8ES7SgiPaW0Rm56Z7UaxmlXd7LTZsixnBz+Sn7CvQHlU5Io3iW9L3FjmPOD6OMbL
yh4mFhQwPoGZDImmuEyy9hpZu3f9B/M+Sy6L6yRY4CZ6MekDUIJNa7BL3otq7Uxj/C17Hs+9iLdB
xq03296FasTQPDDh4b8KIE/zpUWz/W+eoc0uU2HGQPozkQ/38wga+rpKM5iDmTFC2o9XhrVFRR4W
EVEN1nBhiYAwm6UpwTZhlrVidgUBgo9bEka3Q7J+fv/5X+EmKMk+X0cvF6PeWY6bDd2uZ/HwqlfH
jUwJEjuW7UciwEw6si96cuCyanUNDn2nPiNY+USsEmR5RjiHKj07KWcRjzncxI3xTBl6AdfpaADM
stPsJahJlUAXmbGOmaMnYanxvJM4Pn+0QPDEsGgXC4W0UQEzNL2HjCaLh2Y4Rvzh2md9Q4uTwDux
ivMUhC6wCuHtT5M3PUN9Ac8qyAnp0DHeBUo7WTkGgZANszKfFVyfH9NqwfcZ/c0kkyK3YpjfiqX3
+H3si7xR7cLc9KUaox7yTkAGY3rLM+O8EZ0Xrx4fmJOpEppfgnMomYCi/fFOoGtTWutPWJXnSKya
copDzvBacLHEZ4gZtfdV5slhR8N0i3RpEknsQ3V6oWzNdQlK42EMWx7lnvYNRun8D3I15h5NdHHx
INeCU2/9Qmx5+RV34iNF/S8+3xX66viOtlu4iv8Dg6YdXadt8TVYsFwuf7SXXe6iMRCP8ODFPZD4
PhDvfwuanoyuN7VRR0aF7t/JT8RCmodwRbPUjX/EPcQVtF5EtCUfcpskOLTsZx/0D1EeCBZxq3R1
li9MUC2qjhV+naagMkaO/P9uqaK8XsOQkeavXTjfKOC1TWo5e2dXXpic/uNcLGZuSfFJQ5uh3tEO
3jV98IA7QOA9hU80U/mp0QBZh7+hXKzdpRvwQG03cEa6BKgO2IrkhXk6kEXw4cLtIAfgcVuyB2pp
JsMcx2H2T0fzpln/X/0agzjfOdf7XWAQ8ZTRqOd9PRynyeO/LcGIRbdXuVaE+7N1OA2xu/W9mGN+
WrJet1bghXN7CByPSh8cfLYVySXKH2vnCJleLezjvFotY59h1XZ5oNOihyKa0nQFg4Zgmw0FWNiI
6VIPYn4+O2GtlQT7vRcwTfeQH/MAq4eaEkRNuwemYQwMygao8ulAQm/MvUA//QJko5ka6H53eUlV
bw10zQYtwXYnKW1rGnwbamtDEd7FA6aaWQ6YNl9Gn+dmMfpDXtwezWNSYTsUJC/aUlzQXIYMPPtp
eOqEMt6dpvFB0UVKjPHlpF5mUjHJB1E/sYHWt9xnhQFNpnGGiRR+CP/AN5YSnivwupGH2HfgzP4R
f0TU/uC/4chjfz1JPZlEKmIKMRpm36LuMsLCo7KWFwdCiz6Zl9lGBUv3jRnLnn4S1cc6lhcCZMM5
YdZB4SurjPJOq5FScp1+p6KPjVzOCPBrvv+G6Hwu/UcRXOIOE9xmupC1djcegBWxncBDfvhf+5OU
068GVaHZxZ1Mhfw98y4KYP8ORzUSoNIIhFvJP1j1MycpyUiuFFgIeMPPvmQ59rEtC02Sq1w6tiOu
1pXS60j77curFDdZ5lYerzWGmb+repj/BYwiwzNhlmo0998rVNB3s05O3mzBwECCnFrxARzTc7sC
WhnuaizDAAAEqFL0wcf8zlYvZZ8S/Z07TwZjDYcFTRlD648/C8JiRLTslK6DTgxvWYo9nUwtP1LG
GwSM0OU6QmsFHvgh3HnY+1ruiEexwXdlLe/nqT+k3wZZGKnF8EJfJsVmYVr+cDZOt/fweBJcQm9m
tW3Pn26EcbHpArHdUVcqlVd25CtktJcSl0Uqem1ANf55Besiio63hFoO3I9BYHN/Z3DdOSIpfgh6
e42vDNL+U/miFrlM/b8XTqxBjetprIQlqOQgEAf542Wi6EsOl2Gm+cW6qha52xvL8vEj7f0FDea1
SXQCPlg8rqGY5clEeEGC6Czzh6FLgP3xlffxfhiEDgCJNJMn27iI20Xrn1JafkH5Pr6WpjyOcxC1
tfIR3tqduG8pOljZJVeZIdfsOa1cNaeFXXERWC8K3J6/IJ63MapmCI7+XtwR7/Z2d7pYulN34eUS
EfN8wQXJsEbT/8MMKfqaM+V/RX1lh6gWRxw2hLfCvbBw+cSOQ7T682TO6+MpxfsawgD85nduKwbh
0s595F8BIhGZ8AaFa5mdtQ/gwqXpYAQWU28ijwG5wT5nBfGbJ1RAAZDTbGESlP0S7UZwWTEUgdCw
Ukz52GP8UvcBC2PCpe1gXLZHaz7+xnnKdPrDWJEMAjyB4JN4wgUdtBHLVRZOOnYd1vxdHxl4Sb0l
zc7crVXlcmbs/cHLOpz4MaCMdcpaEXiPUbFc1h9thFMm8UhPYEC/7KITWMfCNckVpoVXlpEY7ziM
0aamUJO1Ywf+6vay0CGMcQWbyV6XdlN9jNl2ioIN8YcNJlOFBcKDr16tIRKSBE36/RgIvtspOskt
iKPk9zKsLxfgZEF1KHEk3RW0m8p+boxM7md8qSGm9wnIwrOAHWG0KWRAnRx9amYrGIL9tG+qwWXg
yG44szHSkh7zZgL7oAt7mfsz25CExtqYFBSDCPbHITdkMq0C+pfLrv2+PWTJIdvZzqqyCc1khKe7
BthfLhJJjWhbdfiyzUZv3CCRgyiSY1qpt//0B1vhB5kcjzNuuWvjoSCwCrvDdG0ymvVhXrzbg3pj
UOxuhuZyjRaPGBHRtUh9A6F9Ybe4uRxs4E0gxm84UdQe62DB7APkdZjUwmDWdTBWPdof53gMBxt1
f6hnp1Fsurs16t2ygJOaW+XUUTzbBwke/fgL5AoQwkUScZY7Igy/6x61lYDRXhiJ9jINSkJP3plf
qNYE+mzzgZl+A5waoqbhHOBHTKW++YebXvDFN8dEqMl41um4nyOumpoGvzYWuY29j6JP6yj33ZtE
oiy80kZGpmCtDnuSGJ1/J77dW2Z/ZuVmFHlNN+KNSSigaouI4yHGeUqGbl58BhjM5nVlFNyinv+b
UisuZbPRdpWOc0sJOT93iq9EH+sqZ0lRBNORRHVKft04jKzSP0PIAOZN9aomyF3VoseATXgSPWm6
k4Mw06+uBet5pTpBX5lkFxV+n2eKVfjsg/l3fKveGHjw3Abex6TBPzowT09HiG1AlkIFFualPhNs
tW2RY8oysNGg8ffY8X8G8boTLrFZ62INvdjHxAgFegYm0rdZa9lhmEaPH3uT/rqJTjP7GPw/MUqp
6OxnGGPRD49Y2zOwPXlkFQSDYi1xCouDhuFCc+zgXs+Jx4dCIxhgJZKmeHeTSgPe4EOM367F8itb
RFlnNTVMVBkrTNCgq5It3OLp5mf1TgAKuUZImEMZ/vbNacxcLHWTPK8AvU5J8hLE5IBmjF9YgWhZ
O3AE2ZOGrfC/O6N/nC4NNwSFrecfXwayVUPAktWT9zqNIyC9CpnC+Jy3dVe2IkUy9ISKmO54HCje
y7iPxerPpWiv5tqmDiTVfZbXHe8GEOLO71Nxi+rVslEf7gb1VMjWIYbjA7pMjvNTohIraTv47G+x
gfUrTPus94+OPBHCWaPIeG9CWgepJ7F1mdjCgk59PfMDpb39M6c+PuXgYvGV1geZOHgdvuyjwmfU
zMOiqbW+9jFGaS15Dm1lpzf6zNABfS+mIXwIL20KZMo+eY5p23X/CNHacjHOCdpCUY+Y32oLxtfd
mXgvX7KSjWMc7n2bpM07/C2q1t242jv9UHWyNmu6ZbXWH/zL+8MRTULw7kiAHHmkgno/NTqlmV1r
iO3B0C+WHGAZB9zN6ndsUsieSqwVj7bHGjjyI+t3PQJR6HtwXkHucIyL1h6Yb9LEjuzmiPugVERd
xjrKhiLD3R67+53ruMhRubs1Q42Wgb//N2PBV2inFHr6ZToJIJtV1I+R18U8n5JmqJNrMvw+Amx1
4hkDKuOFqYBNqG9EkbD/isVnEfNkHMfddNZJHqJ1XdxAggb5NUbnniaI0yMLeoLwhpXYRBA4GfAW
YOQ7/PhFZ+fZ47qRdSElVHK3GVAFEf1jVSMtFytDQvQ9wlz6pXFLMFRVtEEv+IEVLHThxC8AN8if
s98wWYHsxTvR+JNynCuFZSly6m7Y+IQWYemWzgJoWOA94evNaKY73h9EvRbeOojzgDS0fxtcp1+E
+6VWTxbiXpTgVgf8C7iTBYSo5TyE7znIcMbdr8d0t9CEdbCHfuF8lJp3Nyqlm+yoAoojwY/FT0Wr
d/cyMTZZN4c5vwPJLHvaThOLz4MiPI7UXAcC0d1w24H5GVVbRBOtMuZmKGCuFv6x6AEWjth/Th/v
U3nMgXN2HAHA6UcxJqHGQkvmMuwC4BODSPb3gy+4S9pqTAgH9GW7dTyEtd7KIFgLXc8d6pa9gWy4
0aSpjYsmktpZ5pUtKo1T/vFzp2zPq1qwa1aKWNzobbwMQtDN5JAqtAHUEMrLjakQIxNC3rns8yWa
Ujkbg8/04O6c3xy4HcVv0UxVuGbjDd9CL2rmCDCV8H6M57pJIZa96xlipA0zeDYLZWB3HQ6NZOxx
6o0ayCt26RVfhw1tJ2V/wpR6lvU2Ymke1ZKxvNGFOYuWdVnDM8Eih+TwcDP4yRTnd2EmIKkZmGdn
nV9xw0bm/FIBHs50aLclvT7if/YinEawbL2vIhvhc8iniMCC63nxQ8P/z3W9wmkefokImMoUvS8V
O5cwtD9Va5uPs7SfgEpiOXu2xFTS/91ScWRQIa3asR9ArIPn3O7HEMdR1ql9/Pbgs43pD/7uZA27
d3DpIhTQOMxE/44IAABa5N04YAC4vSnWFHwOCfc5vf+bxEcW6wvH1e7EuXYBk/CJLvUqJvnAAC6r
ICCZ2vcOq0KJY8F9YrJX85uRdSHSz/8NHiIPcXVxi8GqCYksyTDTvGctMk/AIZQN4tHCz/Ku4TCM
lmC1VLsS8I2R/bYa8HVY/hE0MdtZIh9eWUTc1CnlBbCaosYzQ7qk236pNJRGxAC0LzvE/iyiV0ZJ
WIgGQqvb405/VU7on3Dseqn+xTRVYv05koRLpO7m+h01X7Qz5+iBCSA5Tc7CViCgW3CrnLbIV48O
Kpb+9Rm+TYHC+kEumC6WdJoaE+SiLC9BnrudHQ/jhXXV8fLLldG/wTHOOT+/OTZLchmGUeW662VQ
14g9hbF3PmsbTg9gZ6/vpzdtIIEADRktGCKIR6T3q73IV/gjrBZJT71kq79zw8aEN66nHMw5ex5p
wqz41o0LqaOWEMrSh8hy4EyLNB2knPYw6lKDbiFZFzITQrHNBfC47yP1EyF8ibLp9a3xUFv5WRRA
naEjSxv19QdanHa+/au0qVo+jV3NFvq/+4YnAvKyT1WF/qNkSybD3TnGW7Pru3gDXjOoGnGIlZ8I
iiOrm7Md4KvpYHj1blWP62uYDrA4GjuB9zmrozpoY7zjiruwFUKU2S/q7d7oenvbDhfqGZnRXoly
VfFeEgn3aGwjQLl7zPHgBo/+68WFnoG6CwKeyjVWScBMDqVl2SLESMMnPNOITAKPT+qHnNnFge8n
mkbb1i/N5Jf5qpM+HqJftv8/nY2X/Te8D6eWJbyyGGtAs/Xx8Nabd6vB6wyLcjB0vXj08o3gM/e0
QPoXuC46l4svIJWXMSUo2EizwXxtLXiJFSIRi/UZ2zA/JZMycmF/UFBjjXRKAf0xOsQi+cKDT6HB
3rB3fbmBLhCjTi8C9GAMSzMOHmAs50duCvqg1n9If8NS8Xt5I5YKJC53ADYR1bzeopieDUdVD3xf
PUW1AvCDEGgU9/jyRW4yjqSb/VkZa9gsZunY2ptrkegrq2yZ8A6NfShm8jFQ/xnv+FfqZ2qHE73g
+a7a3/JC/sd6GiZoo2rF6hJhLZu/FlhQEfS7rX+1GAoonudpIUoT83ANKu9MhwHZq7Dh0/oW74wZ
5ccB7h+g+ibD8u5CEqMsnbENWEAXW1s97RNdFh2JSwydc3HEplTfwpU3LJz5K2eM8INqUejJJDhQ
/vRNKXFffjPVIH65+8n2O48yb61ns77uX5k9Lrj5vTMxNWGyY5tO7Vb/IHR/kbyjZz/F4PBuYtRG
4f4sGKHD33H8Wc4q7rwGl4zvZ4OaKsQKELjbm/3q2AmoRYfm2W9AluM4kM9gx8/vOpt/1A+HPUCa
yJW2s3fjQ9Z05jjf72XkzrtzRNpUJuGBXSIO5Mq/JVgoqcb+bg6EcWJj8/9emDcalzya7VBpic6p
R/OeHR9Rw86sbP0K+wok/XHiD5quFnQy2YjzwW6TXpAxYC/AO8ibQH5GcF1zOxcItK4e1u++ebVO
aWRsd3IXzzFJ41cs6hExrOmmJMBNhuSqSJLRIhHDq/34ITnY2LNL+q+J12Gc5m8sczkdAhxwGRqB
gqeNYiUhb3ULde5p16OuF+cuK7dM6YAnUtM6mbzAou5Jk966BCAI6/CCQetAGBxX5twl8ufUQ1Pn
vZzQOibKJ9Gr2PpbQGzd8V2AltZonbH337jfndg32dIMYmCWFdP6nExV0z4sGfDdv10EBoxj7Sy5
5wwxkzLMob1c1kgO9db1F1eThBBNioCWfrOMiWI2LkS7XUY+3sApgPcZbjZqtZTrkOrJll0Dbli9
35ZNmzHhJkMHMhTbBsc72UaiI/cIqm58iifhSUYQdpPjWtAGtj1xqheamQYlZM0EWqre1D3A4+7O
NOFWv9sjM1tFcs6e4/fx3b9mif2IepGZOn2na84oJfDjfl19UhZ1Vni/NVO36dVSZFmtxpvqSjRr
I/ccSGBceV+jguYRiBV71qaRZrhZCNnIaWnyRNyfqlvybcBnt1BcLtqrQ26L4A+mEAO2zrtQFP1A
OKgDTJ0J7nwYv4/0yFTF8WgLUenUjLfBqs4hzZ7w1KwIIvhEQJsfBB0FhycU0QrIWH6fdn798UB1
kSeWym0ACcBJSK126Dqn8y6RzGYmI7ZHxj0teqMns+eSFZUX67fh4yUgZnk4bNQPXSjude14QrKo
sTpEMsVk+XBu2KJ1Zne4tTBEQaK24xsdM2PU8xaOckQzlQfy2zh84I0whFbeXKEhnDHHS2i3GU6S
S9f1rqSGxkENkj+gMIjnu6hbk6mJMNpPHm8W0hiFfhQfAOfKj5UdL3Id8Y+PG2HbbSLfXwZJgY0l
kahkV54EHKm0PLlIFwawdEHeflOScDibj3aYPmNpdMAGskL0t9GvQkhd4p3lUji3UYhXogoxGYfb
xpZ5na9LJPHIz/ZOjtnx5TkWvBZxdv6WF5SrjYAhtv8LdZ1GU8fhu5Bh2ImczS3aMTohUO31Cfuq
+a0n6hbafAFLG0VOjpWgVx3UHzAqu8uqKnOO489bk9OThjzCCGvD3/ogZBw4NQOm5LuM//+jXpKH
0AhmX3wUw+frQsH8B4PWG/ipkL3uqPDYZBZF01OLGiZdqwAqMJRcQDuNUhUsDPovpIP8QSA8OjQR
yb35DVNMSdTVojPMEnGuq77ALaLV0mgbWiFcOBzIKJXgPl+yNuC/s7bSpVnM69aDwql8PsFUtKoa
2sP0mQUaeVjr+l3skgTDzIklJB6btw2kODdLa7GVTJS4PBrWZf9nK4Ch9AkOOgXvFxaw0ljWk8u9
bTMmwejGJs3DCCiA9KofRXVThbQuw3gXyrOBcmkU5NB2Y5Vvq7J8LAXw6BRiFwGFKMt7KmxnIWEx
hEBU7LR8nfa3Sf5EBZV9O1dL1xkkwPs9b5wZ0UH4dxMTjOGVB7MONIpc7xqU3hyNXHCDVFowrJaj
AxVU3FgplbmOBXB4I9IDvxZBOt/4gYA2SCz8h+b1sXZ0Iuy7r1rB55TR92VaBjMc8i0wvxzqf0jI
FxfF5wDQ8W6iGKUBpjg9tLM0S9GE12tNa5aYmFPAfQ4YdaDOXZ/j+X+ybNakxQwPFGv1zFQswKb7
qHGmFuJqpseZGa6jFC9XvpTvK/4NPQQtAg+Z2TNBfBlpEk96jNVTDHc5JhDBb3kj5iD9rUWbaZHW
wQ64zL9rZzS6weeSLIhmIILVQqw6pB53S88vUArCLuZmHLFoGvpTIVWjQ7sSpqseGJoTv7SgdmwV
z8AhAbhPa7OSujDv4FQ8gQNnnqCEb+aLuKpxIlP0/OBZlbBmDqcSAa1y/B/71tiEeJpaXa9zQERG
MtzOynH1wGUqFTWvoAONgh8Z/+TAeyi0/5vukuokFNuWBcwMOw6PXZfwWDL8sKlDlFwB7j+/45i/
EGNwifKPx02qKRiQXGrMaahYo9WIg2R5iPLDXUgPSU+7o/6/yTg60/5NAF1E70KRgTsCR6FbICxs
Kk6KrPN/L+e8bLn3HvRrntF+pERnyrI6YZHZpYP5rHPT93udgoAUv3PO8qXezZI1ZAFLbCI36gRI
LSeZzQa1oVmWm0ccY5ez2NVcDWDXzOss+M3kwkvxXuxnn/dDgR0gLxDtg7pN8j8szDF75Peeh7hZ
pGxKRGhd5Up1BfQaqHIeNVBUuCoqQmmIEEo55gFBMnhexlWpKr3w4I37DV9PBGfHmn/6N9plv8pI
/ecOMY69DFKj3PHqxrIqj3CP/tiZYgoOCqX2Yo8WfoMxlcqJmILpsT2AGEZQTWj/2prcQJdNVJbt
CA2b9LUVGbcffUEb/eggLVO7jxrZAxhfxSQsEoZIHdZ3QWHFSQklM+hJUsZQJt4nWxjw9cMD7XcD
uv06836a+KmxRRAck8zNJEFDrDZguocL9ZlRUXZa0aimKQttUyhCLYpRuNWAu4ACbhJs777/GZXa
MU4CbVVRtyTXveoe127J21BSfTH85CFt9q/7k4hj9erjvucbekTAQ48IieeTnDIUNtks8ZiNJ2JI
lO40RL32DfjIxK4tKCbwv0wJNltxEdonY0/r09/lUyLQc+KN0rQzRCWiHXQLjVUJ5WLieH+BWf1X
KseEqYTpQIDF/S0GSa3BqHrouRUMAl2z8VpqVmiTqVORV8GXQm3SGOcfiWmjRi8v1h8Em2bvrebC
T9iMN67I+EFkBiWmBH2IYNSUZ0CbcJ9EveVK54SPoOCgW/7SvwFlPx4mWgT2AKS7XUAciJUZZfr8
Vd9k/lhrmkSdViAwcgJPaRxRhyu5EGdTOaKtUSteXSdCaUexwCgn0pXEfdicoyHPhENY0E3aheRd
EVWTYSE/FQ9KoKLMx13mtdZqXVRWlY+MfXuL/OXBSThiuj7YVEZ24czG3JgRxWI0QpmBrgu4LdrH
Ywigu6VyyolZJxF6G4UhjFE+noGwPLAxGDkBd9nAZyQyXJzjKDi4AhczcRoRQ/XCGbA3RU9CeKyi
jFbRZUm50YRUqkKXcYed0p4UkbFBFtgaw9zc4emliFptYeWY9nNpODWnhFdMJMjOrYXhE5YbF9PZ
fMcruZ3RJkx8hfcDtU0tBkkBhIO/DqWsnd9tnsSmp1IBxMM91VH916O1Altx6KcnMTq/N3BIk3ey
G5WjBTETNLWzapq7gdSXL4U8zeTTVnaaAfBHW43jVRxjtIq68iaaJ0Ys+kzX/pE7mRGbPxnMKXkF
MqZ3H4hgbpP4d3wgcKuE5L41aMf39BX8SvAHAaQ+Ep8p5Q/4NSVWbAweeqK4J/FyI00km6+W+P1W
lIC1vGP6PCNOQzwLG+UGmzbagk8Ev/hYnZy9nu6unqp+wk6EprgKXX1mhVjiDItybuI940Pcd0kA
Cu5AfUsxYhfOb6W6ycnXe3+q2ljuPZa9/6ZWlmVpaQ7XqbHiui/5WVuQhAgf8JTNNIks0d6f2VWx
Y2fw5eA3WvSIsyfXjYGO2U5WKnW6IFZqBvGcyBKpLlQ/9QK+UfQuZkwS5URIrnjeY5YRx9KkpTUJ
/wjPTr+jIAAVj6cUrN+yV0W++9UOCS42YBVtiyP3/Ft855aXAIsPMJj7b2UklUfO9OeF1Vq81Nwi
48SNGpZr6kq497CiifD35wlYMfC/4GmXxu/fIcK3BIHytChmfgVi5eUmGSjSRHiTAX4F6J6V3dhZ
9Khlqd5acHtpRBwdF18GqlBYOaREkeKwQ/L11aNuA3ekTY2T5zcZth2jiB4zqeWbrq7xOQ5S9Hq0
XpRQ9z5KY9GRbFrBYxCwa0zbaOxx1po1A7uzLGckilzCCc2I3HobvX6tWpQ5j8/3u0wjjmobs3jA
vGf46Wn6LOiGKeC3x8jU67fnOo0XykwBsKGGtvAsKPqXeSRifD/Y0zLdezkHOu8+oJV90n7BjSun
njB0oQ7xR1+CqlkhEFakcppJeY7Q390520beo4FsIQnoS2f2Vw/R45eiRY+zpB0o0FEmo+02EPP4
d4NsKfXBSmBmniZs9KWgji6tHDsXrly1kzkDHgk6Zncrvu2lrkpMPNa0/ypc9CLtANGYHCPr98x4
O/ZWb649kjidOr4Ob5wwiVYp1b/b6izXDxdKomSQsmkNQtFMZdxZ/5DTDpiuCw4ZV7XrvIdr+jdA
3Xfk26GQmXPbtMBYPUQJw/9NXg0BS8lq7Q6wS7PplhZ85sQzWks60WU5uWU2PbW4YeIFJ1MJ1fre
REBQyP6eycwHomRu5GQmF60Ie9cz+bAP9nC9gIXtsHZ7gw7dQhGu4ZpycejudCjdcwYoRcNvnhf7
2j49gcTiFGfnQPr0iYwx/NlJe/gNU6MBf+io6s0YtECXHozdgoN0lwsUaOnHRQPPhqebE8RRDWDv
kue2bc0el7Kst0Mp0GpttaUyxhgynCRVo5jPoQs5fLVcvqHFuKqm1Qc8hRH1aypM2Bm3Fv2HGVzd
cOTktTU26hF66G2Lu3D5ljTEwr7TFnANy5wBN9TdNfNn0S/bNlp/ePB45/JEz6lXFebQLWj94Jpa
IryO9wWzbkYbPX/jDQAJ1ecrXnH7AqvIkOC0ELkER++W2w4f8n8+LWn8qcwQx//cpsnVXxAwyf+2
TwumTSSy4fu6pDQ5XwJaH0wVwdB8QcEO8yWWvmgmS1fsjcr4okx+Iy5avbqI+eoZVAk1Myz9Ogf4
ir1XBnL1mkR71K54oB6+AFBcmriB8NAhPGjidFPnPBm0nwWVxHjtNmfjguj+utbwJY5ja3mmrElm
9G8PYQnEwdGEMAtTBeHQFJMv/rOeURU5MnttcS65VNfg/PV8XB41HuATJ6qyRniQ+JojvSzEdN1N
6gmPBTkyOTm/FhKYbnnNufcVjeMJvqIC8W4sG42kY4dekgukMC54m6qBIXKcMJRvcJ1lB7UJsOtZ
YVr5YCBJltku/SkrXGuWhqfAZh5qRAOrNJzHBO6TYJmR0ay8GuDBVtNETnXwLEeadD067MXqUwcu
t0/fL9WNOU7KHnDh5+cAwdilBWx8pHLGDnbzL/tjhaflXibaoQoDf73S6i5us5MowMRwPztqGiUO
G/nASU1Wu8GUcG+uW2Ii51zvecCL5OAkhZZrRMVrHj7usDis5sxzwDEXjzKYEZRgWUiY39Bxw+bI
EEoB9y5skmyNBSGKwD58CuP4UtcPVS33G4cmjyVsuizxSVL5+hzMHl8zfpC1yvmInJfprFWQ5BxG
t9HVb1GduV+qH21Vqgcq0+BsPiWGmzKRhG45ZX5o41KCAgiEoVaB70rxAK7sJfqnoMPyRvEyOZEH
lXxRoz1qm5EEVRouAIzH2DdSMRQWnuqEBW3YRBS96MaVjQnkSZTxVpV6Copbo3I+FiFfxoAtLXTO
b4aUI2oK/8dcNLhLPcvFhrz5A9bvjHr51J0ut9yAKPJi+utH95PPWivPhMmwD+pgImCf3m6P25Gp
6wM9vofA+1Qg1MuQ2WDRFWd6rB96RiL4n9lLcgvHwqURbvi8CM/iWT9Mdbvxbw3Dh5C0mei0FXnQ
WFKGlvo8zWt60VicPmBS5hEfUejd1oZIA7VKGZEJXxFvZWBH+sqS8s3+Z/mIEHZ+mxxITDaH7TBL
vfC+tUQaLMZjjefRNLANI5iB4ClzRVbgskl6UFX+WjM+v62YRBuh3dgB7WCciUcP/0Q0vT7K7+KL
2LLfcPxzv2SAxd14R/jP8idGV0zeq6VUzqUjHpD28TGVol3Na+KXz6W8pAmW7Ci0AuC5+xNg5GJu
oApdRetlYWta9p5ce7kvn7VtgQrbu1lpgwGzGmN3KvhlIV+MaxaY64C3HLkcP9DQmd43MQAfGzA5
sbqPC+zUjXSZr9eWgwSz+iV5ShByPy6GsVQ0dtDq1JLY2bUXsAPeuzHfJHAWRp71H8bVy8r1H9Gc
b2uhO/1k0cKQll2x8B8jxULLR8HFSIF09jTOP40pI5NfDfv3wwCXm0konbjU6eIkzu2EsjeEZblW
pPQ503FobOT58mV7koxgh7z1TCt1SMN3Xg88yzdqjpRb7o97g8QrWdKn4vOXo4kmRe2ViSZ3dbFN
nd4BKvCyV5LuFvL7IWnpl/d3eMR7Aqx9jKRabTgS1Ydal28y7RdIkz5zv1/qNQyXf8nTQ8dpNEQH
khY431Ez0q5cT7bxkbOTRZPZiT4ZPjAiJqjvvtpBp9gLwNLv2pwnpAzSgmb8oc6KhdvGdG3ivBM6
uN4xNu580Twg5PmnXV/mEFrtDGNfJikhP8fzU5jXogV8ghGb5WHgAJD0IgpAWdTWbtf683nRgT4P
EpaybZdihpSvrZ0tcX03u0FxKHDaGwshk7iX4RyWFbs2/5J9j9AdatVc6a+k5rIcLMNj3/dycUVM
3fo5q8vJfgWDUlCFebN5VB2aAVRNh3GFNuP8LQ8ZAGfExkihDdJLuZxz8i8LDZ+ne56VC2e1S7VL
vuwRAVIf2kbPlHwj00Xdbup/MsEtF1qbsb33KoPjRb+OCChZOHxlGM1tLJk/U30p2WBnndoBDowd
aOVYu9bWo/jBp0mhH3izCL/XvqDDRuseZmAeNuD/D82tXslGwvJiq5ig+rLiOlXsuzAz9Pmx2wbd
I/KrI3Dj//BoxTL53f62+AxSeZolg6na46BjekohyZUJ+powAZrgPC8VBfS6mI76oNR4c7LIJeZT
JH1kCurGKHxdnBF+8PEbqZb67WYBXsx7QAvA8rlUswRp85MhYtqROffdLTAnkzvPajh0k/W3XS0K
Iniy0rBKuzko/rYqlrXJx2xjZsk2aZC5X0np3ArtLtJW9yIo6g5rJXM8bWLR+IRd9GUzKeYVouXC
aq6s5sB/5pAu2vDSnjVnmw9cpC0zGSlHHzaZqPwomOQD14jxQX/wX36zLpIqR7Ai0KqpdgP2qeUU
ofSe/39+Ljv54WM/PEbl/vz5dTSaPyp5KKlXVxLewBkf0gcp5d69v+4nmXgO92hFDHBw3Es3FcJn
oinEYXMlO5rAmmgPLEFLKSvb+O5KbvEmNgBKS7/I68xGb3SeTdcW5vYAoix1N87y6WHjhnE+HH4E
jQm4gVpTCODDn/VBEVjkGR52ASlxfZRlaJHDYJom6/zAA9mfoCbhtL/IlRkB3ojGunvKCVx8fQHM
F6/7te592FR1ZKOgrKbSHvogE9CZAazfVk0fij/R+Ml0SyKcvFcrbbTKEAzm1YF4v0SBLJVlVO3F
uJ3pP5V2Wuvvr0HTl3K38COr0B5190bJXumvnqLlZlxR93J0d63BCJT5oQqKB/tEuI5W9xIuYMf2
4pu0GEspYz3kNQV6INlxuIKf2u/YyceSoHMTWWiXUWjK+9FRahkNtXk9GoETjE5D3bAsgbsq4dlD
DKZ5hdr7gAN0sQmm+e/eIhP47wbuxrcGGrmKK8eTGUCWJd4GyLd4+iluPisWxnziKjTbzo34g/4w
a80ugcIUdCzyGXKXvyQkD8yNOjkqYg/7747J2re6msSfttlGmIewDM8ZLrBLdB9I+U5KYECQ/rF6
XkK+ZuoX/h7wGxUX7dDLJ0Q0acZWobTmYkEzA+1mrezyr2BEEx344qVh/rO+GAOg9ddvSZ+sg9WW
dquB0AfdEN3ateryMT7RVO7S3idCnTs/C9/bv7+juOTjtitshNEu5FDXHebPOgcCIBi+ZoY9KRvl
IPzKS9mclOWVBo+/PEZ8cuxDEJ+0VjeublqW7yEg2mLHGrTSuB+Ze0vxAN86JQ7zPMUA+BU/KBus
tm7x2PXl6w72MtJ9wH0HCSJ2OkT42vlpjgIvPLOWfqulxTlGsYk5lq0lvyZjlvO8qFQKYDcGS4n2
bwD8XiY/tdeyAwiThwUIFos7VbYKK2QLfaiUCmPMZUKSjLwtdIG1CAomeWFglZ9kOyylpS5WxrgF
Jr2FLVwY0xvrDfFcLgvdrwFih+kv8uGcDxi6hqKEU09qWf+uP0esRQ99xVdu+IsxL9MNY6FMjhLX
KgutI3nD+x6+sxnlXzLF3VvWoKCm69sNiL7pIW3CYym25eQ8BKALoptj+AXpGSg0VUBCedBFYnd/
EWgOSxJuFOtA5RmgQ4MoOXDP8FhzlHRPesz0ffaACDqrx2ipQVWBAWj7zyjuOUdkQhjQ6YCJc+yB
b4ZoAzjUuxvt/sBjBfvewfo8ZDuwwXR58InIO/ES+VWaY6bJIhJMWJM9HlrFOQzApZHAqsCLhzhS
q5RTwTKgftnbrADXQDCutqgElRYhrSu0je3VVFVtN7Ef2MxUGQT/jhcTuRFUKObOna4sjH+EMriR
QTGf+CgNSLunpRliszA9MI1yn3v/eQs9D5xDDlugegjUiNWt+G2BPY1xU357DLHm2XJPsCQMxfnv
GuMPn8OjHkKRTMtN9CvMIpBq/MBMeTkHJHexp8dGYxc7admU9bmoEei/1EDisjhcNo87ME6K9/xa
uIckEYGAxS45uRbL6ychrnj3yOut9keshjJV8iEClMmaql8gzCPiSjTuxULPmupucbVPB/dW/FnK
xLws8A+yd02mKB2dhktzCVGmyDwKgbxtAuCV7dqEKIL8sDg0S0mNVZYDyPpTU2zArteBp/oQ5pIe
Eea9vD+6ooavhlmc/B0MyALggIpJUgmlCN/MEFHUw4oQujOVaJz0LC6SqmKrmm2cLUh0yiB7aKvu
a7LFzSujh7OZuMa/bKOuAW2NIXh4CRynrrxoX4vTLl70TeTzjHXgpy6MOfeltc/NCOKBPxOp3hWW
LNEJdEZ4Gw7QfQECFuvl4ABcdDpi7oZHnsE/cwuOZ+p43L+W66ahipA3qHGomtBTRyUJPBCcKtsp
Ey6P931B+xjrrh0jTJY2TUHzG2WhaJMdvkKyHDQplykW/f1stcTVUj4r8rzLUn8QovpV/jA2uIpM
m+YFkraZEHeZHmWevwa9PJJ8KLMZ0ymfh6M3IDdXfDVhUmfQjiv00yXcreV1fnU/1O2UzA0OaL6D
eq2wLvkEh/w+gw1WTI2bP5dwx7DCze5IUmjwgMuByaigBO19yofLD5nQh9RwcKnrG9BICNGr5bCz
MutzDAGpE6eqabaQ3pPPu6rsqQBQw5f79zuKf6JCoZQmqJjKvTzKGm6sGjMmu1V9mzpm2AjnrVQn
RjkHQCQs1vNRjbPPxwYxp1jrUaIxJHiNc7fRxv/Tuyjc4IsMieSMuKyL7FINPzK7GW0IQxBzgNEv
EKWXfjI6pZg/8/FTE02VVsEhMlyAe9Pr5JFsjI9Pzfh9pR/WCppwX6akmU4Lfo4YsNqY5UzsS1ke
k4RQISg3Xl686F318UbHHmUQIGMTo1erLf1X8VnXiWa23t9CwwKgz9+IgM054gHR8mtTChheevrj
b2iRe4PBtV3Gvc+3dHXrAKZhUbsH4C9cWuuJdFBI3WVVBQRTzWOrn9TQN6lXzJ4tF+R/M9+fg7UC
gRetjGdzH4UdQpGkZZ1zuenJE4pjDC0Xo4FH9PrmAq1+1DH+4OdZ/8O/wkbDVMZI5hx6SBtTt5Dz
hikS4Q/4oAxO2IlPhWzYwyaDrKkXEwDDT1Q2jJiwn6kRCTsCHGHybog7hZPvuEW71yEqDQFbFzFe
h4L51qhuiFxp2T1DObPutEtOlcoSZUb8sjiM7Jh0n/v87N2LZpEosqP9oUVyTnR4/hmu09PZjqJe
iyGG08tYc5k18DqFTftaBBRBwfaQKq5yb3G7PQxzQIY7B4Ks+82olXmT7qLO3GfALBmAFFnMvgRp
j/ooFWHL/Vk9NZn//kjP+07WqGHqcwqI3hykWx0wMOU6VZIXgzBGU7HsMSTJcu1Xb+nRXrF1+LlZ
CWn+53dNLVrfIQEQfDDNWgaXcIzsrOplIuv9Wn52qQcpX9oNsuw7+88YJ9ONBGpo4I/+iSpv0YOK
9A9XIObJNhPXb14/vr018he92qd/NmVnQk/14kakmmgAnHqFK2N7x+nhJmJ7k8Zdartg0g9UKYWE
+/CAvuka3I71rTNtZqAtNpUFbxr6AMF4Ed8mBDiRykATO5PuuOasAd6k7y1hL/+ECmRQssZSSFA6
24DOA02t+FyBwJxSqDLYWXrwWmwmUXjGc0hGaymQgwws6mGbidKR0rMf6W/nYiZGI/Gj//QDQLZh
XdvWM2O1uIozI8eVuUri55X2pjtunh+B/u6jzXgpEOFf2xqfdXnp6mwP9guYDXSvF7mJRiewt2Ir
5maRUhDBiRzCYoeqAmZTE7Aoqu1CmdqXBHGBK6FMohHDCeoq69wRty+tFb0fxPiBP6XY+2u1BerZ
nWRx7ZxnSFg+wDFyJZA+jwOqVd8uoh2pKlDt/lutPb7VpvpxYU/75PSIC88hUXzY6JrCdUnMYM+V
+DgMXewYl7njEvy5+BWbC6nJ6tytbIk53W11czoZGiyFnqFFcyzfXNKyLsujlFSHDSnD9h5zl3Bw
8WUO8mS1FhA4NUr8p86gywJpbt7xoxo7HzlHL7L1n59sKY/2DUjbWKFInrHkC1spR1uRf032p2xJ
qIuZtPdXznOk0XbRd9/arXjxhkriL/PEWKTQQthwIS9B1Kf1W5eTXLCI7XCJRY8epjz4eKySOtDY
B1P3kEc14wXUdy5Cvs/+q4s9Zl3gIaDYu4TmTvWzi3EsdID3T6zXNY3yQKHKU6AFbCVvndAEAICA
pZcXWAHnC3gcD40U2e4FtO+FzCXB5PB3KNy7S8pZjbu9RkZIex5C5LQx/blEDKH1S3IeD/iL24aA
vbj4Q6tHse2VK5vkcXV4eIWmbV4XSsQ3soDi4TS8i7L1E9/n8DpiMt0DvQ2EFGl0pyafomT3uSbj
1fOMR0CAVYHBbCZB3cxHsZFEmhYavlXCpK8vzhyAnQH6COHnYtO4VLPv2HG0uqPXIT2et2cubURT
SeN2wu5lLD3kRW5+Je45G9CYOb78WVYFWeraoEmL0DGEWaPDkO6kOwhuDTP64KPtlT0QxWVXMp7O
hWfMOa9yeC1k3NnMAA/hQ8g3UxJuVfTQQFN1okGuehvPteeY5B2BVzkbMNHDnApobkKKSs8Se8vt
kTyHfGp29rtlyiX8GXlKOo+TtStkv5zNqZZY50T0z21faJ+BTuzliQ58lpe4RyStBj3Ud/QU+9Sc
pM5xKeQTJj8usl9fWXcxKGE4G5ytgGMLJmwhiIPK+NLzPLppIIYNEULEWFGP1ISvfZkdDX6F5qyB
kItppi6gXxEgya0Z2pK5M+49iQA/yo9G/DgX08WuLREI+M4czEGGrcwacvEgQNbacU9//NJippVH
ulVBnlO6TqOxvbGC1eef8Yh+4/xXLPx51tjwAHx4suyu1bl+4NUJyWrHFQ6nlCjYwnMipwPMiUXS
voDeeAaU/PFH6Og5fj5AHFyjdUSyTkrLzk3/pbTzbP8uKuyjff02HZlL47/bL28UCvnzBIi5pMNK
hVXfaEY2F9O/HAJsrBRQnXs78Nmr6Mk6Dm5mxsgJGHbolNDceDmHZYv/UANTcw8EEhApw9i2YR+z
0JffPbCc4hf+tcU0GWTczfxJ+Z8JaJ6d9eqCj2B6Onz+RLawbuuXT86jo2/6hsxFzsY9Q68xb8zs
64FaI/J9QqWJkawM+vzEAR5kx/oMfy85FmlEtut+68IfWDPfZ4xETeQXH7PwWqfW2e75YUPL9GJh
ETURtRQWNJ6FXKZUkRqgEWO/WMLJuHS/Lh2aMkifYKJ9rQ7p9ad85CVgR77P3XXGT+lxr0MO4rJw
eeI8gKJ6V5tGH39jSCWlvt58ccwR5hpZLvlACTQlnGuZFIYg1Pf8EBZ0m15I4vZwUHh5hvt/KZo1
AVFBZPwBdnTfxxjWa1MDPf23v33XG5kbfw2Ldt/p5zsWNVf6E/dASN3nlja7aHAC7zmnb72dsLZ3
tO6y0/ThWIFviV+E+90UViWfRJCDY3gTXXpgp+SvFd53GNLg/fe949yCV+jJ9WBmDbYNZyjYc0Yx
g8aJFgY+PIbi2a3RpMOXiWhkryHrNucDJ3RLEujLR8ZsOiaJMwcACw2v9hU9lnVkxQu0LcGI97Ws
aLDMwnhaH4byNNBeel+1cZs9eprf/H6+JcR8KZ1Tn4G7TC898TCOnfFMzdyPpF4nNXHi53sMX/ax
WsyxVOYlAT/J2EzXcoN9cMm70N4ca/n02FQh1SCTb7DFISFoHQEP5CuTRqn1zyW6BGUVqcXKxlUB
MT4//RtAoVve2EomADh8y7rz+N6pTZtsO3iwRsKeR2mXIdwxD1K+aBPvwKmM0BKGyKUJf6aZIWAF
urrNPEMow5nN9DQp/TrMBkBr2t6GAbIwuoPXamO/yms3ZrbnCSoijpA/j09FjpoKq/BTptdcAQQO
vr3u0QcZLh/+Wl7wiCY415PSSesEk5F+/2XF1qKfzEnNhCw0N/GZnnZwHz7a1mfybzBcnYgFMQ54
h9do92vtATjQhQ8rD0KVuLx9rPx9pY5/IKM3cvbyZznLZiDdTSaoNSfpx/+AbZKC2j31VwMFAiHg
bXTa0KDynKMebOba0P/TmlrLa4uv6qNRmQKAKmcvxVT7Dd2vMXVOO1eJuhaxZY8lOxI0y45ZFlHj
PPJsWN26NFWRTLsGLHbqEy60w4PccYIOqFO33OapVUS4zqnpBxOLQiZ7Ya7nTKq2F6i05kV1O0GQ
h0z7JAeg+IFTmKB+bRVWESyg5e4PwUmtzybbkNo/ip1W7awA8mAjj5mCyP6ljhwlNIt4VurSOiNK
fF3r0UzvUlTydPbH11g8GeJXxHy3eMevb9JVB6B57xlmchQs1QxF5u6mqVtiLxtCiscWdCYCQVB1
gtkHaofyUaiLL4NV/KrB8dd685Et3GeGc1HSTkAFkjKahj8TwTwX935b1zS84IhD15ET39ywzo76
uQ4/SLKc6NS65KnmC2NtZMW1rD/sr/xNxekTqiy7BOAHBjygTzGsoXYVmFxbZ6+sHKWfEcPqgpfX
zwDTWfICAH/+0gIKiLuBehXUuUKT61tL61mMKKL2+5hvI+fypGgw3BROQr87g924z728OQkT1p/U
rBsLUUgUBOfZAAbYd++zXaxzXGFhe5WgZWaOE75b0oMZzV21M1Z5+XtxQJ2nbzlekuyzgesl/Q/K
HkhukHwn4WoPL8zMLOu8ZD+yjULEnuN/Y8Ib0j4cB6SR/N1QvlAeTn/Mn/6DAmHLJ44xYvWYsOBi
yaPEqD2s34GBRzA0Ti0XTnGnGXsGAcVO+B+NeJBQHN41blcX8xVXoQAuBMi9/azwFn+sjRLzQLPm
Ze3PnJf0+Jy1J/YwQEQgqvMDpp2o1k6CDDP1tatAAkjCDC/aeF0/BWkm1LgkbBGcSZiM0MZbhkTz
O24/CaEFIjZN5tKO05fCBsWGGid8luRA4z3uNow/K45FtqOgPVQKxYEA8fpFppElxUSBjeeY0AgZ
KwOUjxFbbp0c65A7rYWDufCAtJ6MC/v8HmVClN7gCjVAno9Nav1Kk70hBJAOy86LGfTAZA8O1TF1
Q7HqEFiCRo0P9hl7r+cdDfdT6fL0JEbFz2o/AMrhFASz/AVszYzkvB6kD73Ney1TrnA+eQx8IDHd
U4XMv7VqdywGGEnaLFPJhahM4flsTbyUpVzvlSLbrwbzmlHHI15Dsn79oSgchksgf2wTW/RA0xH/
k/ZEXdlCXAVeExT/uqaN51BCp+YOBvtIKQzBGqA3VabQD2TmirELuS7NqiYiTtIccY+X+rNWzdDC
sYpNcdGGE6NRwcYKxxTkeARBSK8fiSef3JvIgh/eb2IKMUH/+rCHgZJsWI0U2O0KXIgRELeOYLwh
6WSM6QshvOHvtCMh2NnwIOD7xzOj+5eMZ7YA3rXrNvkmMZx8eRNF8xz4ENjQuQh2lF+M0KitH7vs
QZ9KjiLtpexVvLYhaVyiazbCV4teQxc/UzLgEf474AbRPJx1KsIiUkBDBowit2pqqXsiD+0lFoZz
bAzMAPZzC6Z3SpjqYeyTkwHfNlXsnPwnYEU4Vvk4IYfTKjxJj/l4TPzQ578MYvS7lanniPGFVsgo
KwTncPm/we8Y0nOuApn7laECJd+1NZmY0xBJGfYOVP0xnPwnficfHBvNoCI8crav8yYCCXxyhjh2
kHm/GKHlNmALVh3JXQV+7efxm+g+EN/QxdToGDVq8pny7S8BMbDFj73rJpUia5DcSfm+TscgKwMC
Oqg4zhcNKP7ibmGhKYuEB7b0GAp0GSla22A+OXxTsERenGSAwThh5J0xNghaV+CnuJOJGTWwOeYN
qv+rzX3arMwgofkRaEJi5yJQfVdOPOBTIPmYCpOaGtVLMsAqDtrwy3djEzUe8yvGuEF2oLUuNceT
/rP/BGC61rFvezxxGf3rBZnToo8qLbB+S6zRBFvx6ZaSUK+b3FAOennIsGhk88ZS8ESZzQA+L+6n
kL6qcZ6su7WJBKZVWDZ3u0ru8ylqqJkGmFxHP7FDCg8kOLAq4UycduxBhlDHsQp3kKWChjbvOM3H
w72/WE4lXe41Ens7pSMzHLhtXSPNX29aDx0fasVMvtCmti+kdxXzHbtu070h161k+kbEJYijRlBU
f+i5hMY5+Ij4tVFhd7B4k2rzc9s7DJ7hDntpWcp31STtP8YineaRpY/LgC3wgg11K4gk584RFwcM
qxcM0c4t60GwzLzWJn2eA4R8dHJQBIGHZFn2MgWyLpOFrgmXInIg6/r0XJENSGcljE4N+PVYmc0N
4/hBlVW0dipIto3XioE+3YEIYg+ZUoAy8NLsjghWHf7OoFM6qhlZeDU1E3cydK+1mMWUycV/QEia
Kl7f7OZGGzk02iMMjH0pwV26aET/LOyIrWbnAkQMhgOCc/mnzEs/No5eX8RUzdDsyu51gD9LSbXd
v7HsJWI8SxVfZyk7feFfbqTRnxQ2j4gaAYA8vpEQv0MnU+UbIXnHRL5aBexCsOhh69zkx4Pfm65D
4vBFc1Wx+UjNZateqg5htO4QHCj+gEgStQrgrSioTky4Q9fbAcE4TMVobFrX6jI70xl1TZXwa5He
FLpbMx+Gvws4np4gzjOTMqeMVjHMef1iBDq2GAn/4b7WoeMczJYpdwgMwpEoVnKWBGOf+UnpU1po
SQgNCToZEhci2ZisUKYdUYvtNSFqxegCkmPpgOidSg2iqWo0xj7NWFW0i7kLZu0/ECkxmgMiGSeA
QoXorBzXJLWXfZlKBYFHdG9LrA4hK1R8iR0wQg6M9VqCH4w6A5juLB3G3FREgy5SwxO6yNm21uCj
xxBEXz7y60oKbkOPwB2A2dGbl4yhu1qF9oNjG71WY8D87qHGT4xKCXZv900PSmX55BXQoKqNk4ec
YOu+jYtaAd+YqdnR6sRW15hkeqqEq4RdoMFEKP1tEDxiBpONRinEvkahaSrsFVgeCf/UuPuJeX8U
kh+qyy9Wr16BAxrUWuQ5ZpEkGk6ZmIv5q1oUlLbmQVTBOOMjo9tJA+XeqGZ6ddOZJi7xzqkb0k6k
N29iNP9KVhxFxuOGmhvheJ6/orWQQCSsUoyeQdDwTNE/m4dB7IBzzWWKpZyibH49cK6jHpYyYo6S
l+1awEC1e2kzYvSazxNlRJjIubzchHgoJvuR/kDORYFD3BMqGEjoPx5tjIGY7CsqWA9L0doBggpf
K+MH8WaDjgLGbrccXVDgG5sPTy5r6IXSXHVgpvxWERQ7tWVmHRti+Oo9+6gMki73T1RpnUiMyj5r
RaI8AvXkJnJISCwGmmQnxcGpHJMz8jTOtRfIaBHpcQJxfLwbiHJZgitK792eC3u+hJGhuj1aekHZ
p5q/pQARB+LcNiQ7xr95MvDr0GgAyxgjVxYYWCs2X7X4wPB/oSa6xxd9uRxjQ1nFm8vdQhP6sHIm
HTT03PT0kuR/G/JPpfCw2A/F7Z+FwTfLCRLhn+UHor+0xjBtGhKRTF7XX77Szz2U0B3BEnuiZ3IH
+zEa0kLruSH+9GFuPkW0iJi/QPq/IbwlZ/qKGD3vksjoaWIs3bz4HgqeLCdC5BamkBWP4Ei4IQhk
Oe/tfAA9Vchu2LBIn/VbFFXsVrFliqmbJAoVB4GpAaWeLwHdZvml8mPYfy8jvJtYk+577vNQmSzF
uJQq0x8DKRpyqNiauR1Lc6HR3WFtehaeDoAEDtuxsCahFO+nLQvHrQZw1q47gYFpu1Hl6MLzkNve
S7ls0ssNGorT63BkL1CLJkzMnHy9Fju1eHtD14uSzuO2zbZ5W9W8RSlSi/iDwqngGODOA+tmzPht
Z697RDltpLH2/zzlkIxCE3ad9vEq04wrQTfErT4mURJpzigL/gLzAHQqq64lPUXGtfcdliXIwVbf
eokSLU/RlJDBSYRtIVKAMbz5PjYyn+yAUV+QZ0Qt4skGMppA2PxhhX9UeIvG44NzAdy7kbFx3gpj
KKEnXnrgZYR3bc4JCaAu+WWWboB9INPnf+yiQZTgr6g3kUEt7sbLTsNah/OzDbPreRnd3EgaTUyq
QcqLjouVYTGEpeSxXH7KQhIizc1iBntAptYNHk6SAHnE+W0CcVNCWRwtGNzYaHXSQxabiSxyFF2e
/WDTuv3ER7Wp/gI06Q5Bu0wlav9Y1Hu5vnY00xcqAwhUIKTcTmfbwh5vEyiaepUI3VDbdr1NAYWp
DmRtsJ2wFaz89XcaSrmeO1qovOZEt6XBLAbXP5h1X+u1jL8psNLiYFcuOKRR54R/iiJmPKrgnpJK
CGFHceZDUlaqTbxMq4USpfoxWt9LpAaeDdZG93ujUtdWE34M5dF2HOVkHejslWf9eTHkSwOKMCM1
PJBZz3hq27USzlNEPTeaPQc6xN9cMuRVeNCumf5IXy2K5xm+PfeEva4iIB3tDbfjkghYP7NTN491
JuPH/qkBIl07HvegY8vp3BMrVIi8pknYU40XerDANJxhB5HWXy/mXgGQ2NCf24S03tgJYBjBGyU4
S16aMM7IyJzF0ITv/j18G1esFLYG7IZ8ngK4Mjteu3lfdclVnJn1mbxTdelJsfVZJNB6Rn/9nyJo
OOAWzvEqLZwme29+gIGXe0waf+A9rpSwU2npzot8uUeJmWG1hOfJ5492ttuQaXZSlPhherzBLN7a
k0eTPi2AUaX3dphQY2ligoAuyhi9Xgiy4sQCG3YBK+HbQJzxad1TNuBFB2R734yvKlcJ2jBMwjZC
ZF2O91c+uoIQGX/Hdsgk8ePQ4VuACE1MHtudtuB5aUGTnyEdQR1WvDKqaa6WoG2PrRh9IB4WWj/3
3ZyaebM+pDm00mwnqq1YkM0UpmKrvbowDA/kUqR9RiMH2dZ7l7iXO0W8cBY+0CxmwXgeubDTlTwZ
5Sax5CVoDUrBQcNM9go0MwSr8L3/tiH2DBS5uBMgEmENGWFRfQrRVmM6dpLjSjF5YSYr3K5xl83a
zLv3NZsnU6TRvWHlin6AylK3SItirf1S5uImlYRRwWjcyge6Z7nZjIEHwp8WciumcqvoTVfgPA0g
5k0WmUHihyOP8p47NpLnGgmB7MpM7CI0VwQig9z42yQJEP5mr22g+D5GtjFpk9bh+0Gp+nhxw7rb
lnfc1a1GewBbO+uZyWtZB0nKENRcE4fFYAbK2G0Kn9e9j4iQENYkYPCQGTy1ghZFwFNa+q4OVfVe
eQ8xgHTGAf8opnZ/MtSZniTgSstArLiIGCsj4qOJn9WKreq6HKO5647sViW+RZrR0lvfG+9BsqeX
flAbKxwQSUrDgBg6UynKqKEcb4j1ScfztIakOci9rdj7I0ZFSdTeKdhA5/DyfNZ4mRWo6f0OQCQ5
MmxrkfCYfmLzsILEnrKI01j1WEIbrEUVR5ypPlzE//aQdfl7OYYi00L4bWpqSB6bw+W+FHZqxNoM
nxQ1Jlg/edAZsJWxhpatoWd1C/9dZQW5z8qMrMWvyb9xLtq+5W5e7EK+ama2NMup+uGq4vXtnEPs
Dp4VdorddP3z0Wb2J1RYufEJ6M1MKWR5Io7HU6/aXgPq8CbpSMeDlN7eZ6OYULg1VphlqyqjOF+b
Y2TW/2PDJ25JkNlmFkuWlh+Rf7n/icFSff14L6sk97zeXa/TTXSoHYxG90BbitpSOORINxG9kRle
6XR7vJsUrCuYbkS30M2Ph1ZK+OgZfbB5OQSce+zEaGzNH79gW9qcuQEflAsjSi07Z9TSd8om/b0b
nHg3EAAgVZ/l6A6gFZ+m1YEd9mRqULrzPrduuBzcMH1DYmMXtWqApsC36CzFU8L3AihPetMlDQLT
6BaLosQv5No8Q86n10trdareMw49P1QTp/zsc4Zxwzgb2uasY8+i2kyzI5mvZ9TFJuHdeWik9br2
vnFQ8svKESYzzu0TR86hHxBEtCk6F2yrDke1y6QPyM7pZWF/G++B698jDg5jq3wyyrXdSPv+zoMO
8bOECJ9+AtOmVprF65gqEITpuSRlBcoH1b3UxzDkMB3iLR+Q3WNOyJulb82meOXgZzUDSvi/iY+4
jUPe7As0acpeHSv21s8eLv4W/8PcTGMKqS8KwflWnaqa197Qmva7p6FgZMxt8fpGNViIp3XiCxqp
ml1E8RgxbU1gB/P/ofY6AJG82s2UTtO4JS3PyiVaE0669P1Foy5/q9Q8HVxCWJxvwRv0/wwg1ZT3
y5Adg/CDI+Fe5j9vvN+R2BnW3uksguRPwCPEA3wcc/kEl7pErdLHcGzqEF6oOUs6o3xEQnYY6Rxo
VGKsUWYkTBZhklzEw1j26GeY+LCcFIwi2lGyRmF62ZlcX069gQWhDBn65YTEz1Bg3B3L3mQqmm8x
mUngJq67ngGJdt+LPLaJe6+tIkepEJzgWIegVRKVqagFbPaSRzpXXgl05J2Ldfyc04P/KiV+Y3Yn
ctj+xwbamu5ff/KnQ3zriulMZhDDtz+24qea9plCfyE2+JOUYF2sGkOzWSrW5GT8CtZo4RG77uJs
ReYp29zErQ21ThnrG3AgBDbwJiU217uDTMsJnVQikmHwwr88A7PcW8pMEiO7UY5kSbCDZvpztDQz
Fk/1cGas4O6XjNYBPtL8p8jubVw6AcFsmW3vWgy2TfeuqL4tnwJCjrIPnGi8qlZzAu7TMOu9VDDA
zizmIYzX7g+ea2HNpPmQVG8Yvk4K0hmz5TrdAto1Y4urHrVxMMfzKoj1M7GPPysc84B8svB8CkXw
SNuFKMJCQfINpuUINVf9MX1MRSATMDmKW2f9bE4q8LtG2JziEYQ//NMXwsqDuVznu3cpYGBUq5Cs
Yzm1NmfMKwO/JVYXXOYFLhkYNvROd7d8NJZHV9M3cUqanCsAcdEFLSOQceNKNzZRz/DcMGnu9zew
HYBezIt83/OfPW6+ReiDydo2S2d/isuj08qLLoQttEEnHATwgAfzkeC71LYg0IEH2Age4mb67l0V
+EHn0CTQfdg/sOZMB0AleEBWuCPEYowGFfKi39baHqufBsqnfsJE9UmwaBeAqXxoiDjhnYlk2MMv
hDKQ0dHILlaZq/32D70+F2J+GYfnSQ3dvzx8+J4kAmk3dHux95REP7YMmgC74uRtwTNpSzLuDoRl
+rJlg4ToaUqCN2LP1QokspunO7h3cE+d0gItILLjA8gdiERI7mGdMohzx/lRX9nPvw2r9qt+vIhp
pW6mc2RvFJ60QDBpJxAqhzzOKPy09epOuHnSisbK5wLZn10FvYluRqrMIDecS8Kjcj0fTHOI4J+r
9pjS7N6vS717qRBkfbjDHiKo1DyJe7+W2rVTIhS+NwIojQ6h/B8YwJ/Cv7ZTYcW7TMzXh4ak3v0S
FBwxHtPp4OC6L3hCqUL5lLCIg24KRYftrlX1I96tcb6qaWKLcrlihkrfZpwxjxICQRnuKW+w3psM
RNtrUsizUI2sc+RuqsRdahKklQa7WYG64w0a511NDbYQ9Wlzj3ZXvvlAy4ieWsxRcoU5oi8LQbsb
iekVZMwkqpRoA9H18LALvX3u0Iv4ufx9uLch6Tsfgn3u9A2DLso/lGSgfe1SRZ91INC7pgECIXLD
DVhMa7kGciXpKUjdodRaRQ/9GgEjd+SHOrqaigqHOwQLb1DAieq5giR8kET5bhgnLa9Pi3XEV7Ag
pE7QsDXhySmCZK4Zle9WFYNDEcKSmj+/n/hRJEm1YbmZ2Th9cnXtY0yn5s/XB80REmYc3ugmwDfx
OQ9Rm6LkWbLZrdAe66OsQo2GRxjNC1P8hbOvHAoOjjMxTiEaoTSz14qTMI5VSl/y7M/Ba/4A4QqP
ghSqwVdc2xhAgxDuPDbH7NyyLR/4ZQT6bjaql7uspqNnDEn2U0U3M1i/1bZqZQMm6c4SvhcDweqd
6aJs9K71b/9c1ld4L91RMu0rH6oEqmHHaItWcSulUsg8fgUS7T5SFNpzvMcqGT7Dx8gufu3n711u
bFxDuIMBHdvbd8TkMDi3+AaEbeX4ImXD8GPYufqpYR5dgJ/XaAX+sNme0g1Os5mgFD+PrMbDmkOO
TqNyI4HKqitF3yDvkVkw1kDgbn3tihABQVQ/oTHhXLZ5zj2txE3BGeGrlJ/1x4U2Gtqzfcixh1ia
Sdo8e4lF2ng/m9ulatywbao9okiAfh4K/YeUOsa84F+NKw8v3MEly2bC03ksLiEpntX8Pc4lw3mZ
roEuN3nc1sWQBBTGFtIjr6IYAdE1+cSkd/6ztfa/eNsDpYpntnTPEXHd4lDhUAMSFgzRI87+aIyi
1xokNxYz1ykf+qyb+naCO2JXxkmZ2NdTXfQHDdRXjSQkFOUYlLRqGg0yRcEaYQDLc8altaDAMVrW
wb8MPIiLE+hKPijnOZxMDIICE9+GiMRdM56pXipZOWxlLWiuNWj6xw1kTGzhtHKy0KdHxXyAi04A
6cbVqUo58X5e466PjXs1pBPFz61ti2bS8sVpM2/NND19UEXYDB2OD42ldj3JGWUEK6FWAhOrhNps
Zk2LFzj4o+ArVeMSzCOl16c5+hHyMX/yhAC12W0avi6PGnzAJ6LBz0Z2Oyp37F7gtLlYCGj3tnBw
IkDKlCYGCz/z7fUVKbt4C2fjjCOKUheBjIPf92qYh9IlC40jTr716eFn3261T6estQG9IomF8PiM
1VxohYDflZghtEjSvT+tzrZ2S3qARrNMmoVTAHbljB1OhAwWw77nOGSiASlO1VLS3gpWL1TdXx+d
JxKDuMY1ddjZTMCEUd2cZl0VojIDmey1bvZeo1rTQDz3UnOkjpzDm/FIc5dg1M7XFRdvfZwypEPd
0eFH1xyrJvgZus4WA6sbshX9M+XkfK1yx0uKDux/wO/Gf3x5WpSRPLgx/Qkz8rj9JJ5RkUYO5IIA
ghEzL3le+YPLZhmWiRbMAScFKQajhWZ9+aJHVepxUJDKHwcrFBRZAhIprXHGVVCY5RtdDpKmo/Xx
WEPcwcxLB7URfpqynq5D/o4Ga/dp/YMCfY4L7Z86+xWd1xW7/pQ59ksZT7sYJZv22UmsMjutIWIN
BlRP5YIou2kbf2MsbPZhYT8EQlO+Y0CToTLLgbRk5f3khlAbRjJcJXfySdw6J/GwJbrVO6wwhQ64
uLvAJAaJqfn6IxhpH2jAnT9fqoxdueHXpBrdEvHBPMXSzU58304BMuB37jQQIJU9BkQIANQMtMIB
buCE3PF6kPF4SUvcBMOKr+X926hZkB4E7A8gHJe7L/SZsP8AEjGSPA2QKUDDSapQ9UCm/px9W94+
zmwjQgSiIrKv2WFxOEzaepm4Colc9edKye5Y/k3KDMrkaCjyQ4/myWAiEDNVS23RLPSExxccp20Z
MPBlvfukib/fcclBiomEcXgYa98u7D7QH4n1g1mfc1WZR4c3zml/lIHdYtde5OrG3Jap6vg2Hp9m
GG35V8jNTKR/d+2c9jilOqiwiflLTP8I/OlkL08sM914CDq/5b67nTZXn9GyMEZeQnmBi6cZo62G
zyNooi8wn53ReMbfpiHPn/zGU2w6UET5DRFSGFkA0HLV8k4J8yNOa8qJsvIXmu50q/mLzbv8481h
i6M24G8LZPnBZriak9aMaP42+8dn6IaIJQA+g+/bpmaYpBBOf+oO3mcd6qhU41y2XbGFSfQyFRjk
ll4cazFA9FgA6de0JquLNPTAlU5nuvd5d7cy3nUF5tlvFO1qJI3470Qbi6P+WKpff+f/zjEtMYWx
ElAJN6A+vL7eirFmc04V/ZX2KFxofgl67C8nP39VD6V+Gf23IJM1HsgfHJSy7GbExH4vkVaaRf1E
AJcxAvg5ikNNWrHIVf8svdaTeXPEybWyMNipYzwTItnUJBnOqnAV1m8IpeWSh/5oeoSTTfTTuI9U
XJR1PbOsqT39k8Q20qIPqQ6CuT3mHLd+hiWYJKGgkV8r26N1CRnrPtc6eREKouF9r7wOG8Yf2N7i
bCtMJFC9HfHhic4IB5hAxufRBbxsGjAdvT/c1PfilXor9q5RLiEK9yiPSICz1x1zYm87unz+ZDUB
pnCsDpNePIHWGdOoei30p5AWg6/ydogGPOwOs25RhHpczbLiNTMWE9Wbk+fosPbtwPnWGNC5B3Zo
FjaXUcOHDc5sCiXx1z2YwqovlPJmWkPAlZALEVPNot/1F6gglmVGQG0oRYGW/DLOpXbwHub5QJ7o
GcHNF5TwpLzNkUlbJ+Fcjt4z8NYxOYwN37Gbit619pKtbiFJ3jJ+dXPfvc+RzSnvFgD46ln/uWF0
qhfZLnU0NtQuT1EcKItksW0T2gSPiPuK+l4r9WXm7phUt757ktzndGliSNiPDzqSxlvk8xb7C0DW
fJRodE+JrIeCcnZ6PlsGFA2VXb1LM8Ili8zMJwDcsA+XUMUpj2o6Hlo0pCTHa3Uah589Y0Q3vNnj
Gq+EBXo+n0B+60pUK77BVoUqGeiR76NctZfmfj+ucDmhk5/+NviYLSs2Bq57ikcAIjkFjvxYTY+V
ekZodd7ZxHKe/TTzxwPNs8z/XbHIB4HBZ6vUBwMmQRRe/4vX7UNQx3064yPaQQLQnRJcCq+Hlv4U
qyUTV90wRlsVMgVAz/JZCOSoTQOKpsKnoaMjseVIeKA6kyI/HpRFEUImAfYpovO7ACVsf1gCQPSG
jsVUxhGSGspWYXEfVdB6dTXH3DvLZjbHFUYozXDHL6S9UvDB9qB9QqiG7uO2XFViySHWcI64587M
DysDQH3frJ8LoLXNZ9D9oqW39Z2/JO9qBqEgjKv9tm3ILojLgA3NO2DB+XtlOU47onLalqyYv217
kEC5m0DJX5N8SGvV07/u7drqSKNgoejXbmE2TQTJ3wC07+g6/pC9CsXwqIylJ1wkDErf9zxDxww7
okrS49aVYejvLHkj+1FAeI5EXa2uYQyk+GX3oXAA3il5JRveDrDf7hG66myzXAnv9ybXMM8dw0mB
lwQuCMFU3v+sck8BDum7popSd7gg1MRafpeU4UcoqI+NdFgZFfi3G5d3ECdyHET+cmXFBwQmYtrV
WxxqHK+DhFOYwGQJ9pPyO4CHZOGmNFWw/7ptO0NfqtZRqB8GhG6yXSG183ZSUwTAAm0L4Tfpnbl/
qrIz0o0sWDk8sfBgh1cPy1L7gZM1hz7KgTeQ791MUkuo/XSuro7AMai98M1hHfJ1xm5rC21vSLz3
vgt7OuTxMhmXqRbiG4eFh/q8LG4GIicHZZ1m4UgoOz0ss7qDgf5LQf6Bj4y9sg72wmZFiJqRVNSu
450OgVGFbpfWPY5RvkAKv88IWoL6xYW+skTJeqXxfCEiw2PStjiRIqvfluGK48yxsV9Y5+erJhQl
57K6vJRv5mW1qtya9PaccSCyymF2JJEbYpb6k24gcN8IBn9uAsmN9uJtvOIeMqxMbUR5Ki/vr9NH
rk0ZlgUPTtnsw3OyzpjBgXwK9NzOWfcbpyjTKvPXcXxi4fVa4Qn46jEEtmJzcct937GROOum6Pm8
nX6BqP3DUvNUT1rKDZL8b0+S0poqpoxxhaz6psUmd1/3h6x7Bex+6fe9cibitX9hjwiVJ5a21d/C
jAG4on9kXHfADLCHiXoxbkDCo3TSJuoQOHp6k/FIJ6d4cJDY4A49z33bvdNCmgn7+nity8JAkuQo
k/4/IOrPPFb705yuboKCtMqSLxAH/SwR3Mrq5N16O2q69RoC+7AVpAbY5evQ0wakFotsU+ZTw6hk
LrUtZXczGoZeMtwVu1q9jmWko9Kw46ARtUrq/tiLDfRU87/e+/wF5fQkqLvcT2DDz3yFhUoGNgyw
lZi/HSsYGGAn6W8ixSrqJaj8pptHvp6mq66O84kWxYTZV2Dc4HW7vThuJ/heGUcrPyesGDSCdqDb
foYFLcIL5UpT6WGZqkGFDjwfw9Hn8Ygabyc8IGJGuC9EhT2oO44LH3ikHUgV97w8Ks8P2NdfK88W
jxEzJ5sx0DmqqAOHTzbxZCFaakxJ+dcH33c1Fj+PUJqMXNlQuP2DYLNjH0WZ80pqxuyPubbuJtWK
n4QzzPxVYwyWlziCGhk0fvr+KgcZNji8mJygcjA0LuRZBN4hrqS2mn3X3D+RzJKsPgFhRT5r/IZb
Yg8b9R61wFRnAXkeVpSge0uKFw7gZJ3M9ruATk+ky53NCD8ehsaYB9XzvouO27AHeKnuGuGOIiKg
4fhy++6Tb85ipOr8wHcwSM0ZogQGtAipCCMYlQcfZkH9pLcy7/dygdco7Q8T1Q1KRKcvjyJmfGZs
gvet9oTqgehtSTHiro5tWYzWiqQCJSeCocpfCb9rZlCg71HFXmg74rIdEdqTxil6r5cGI9bFZnr3
D6B2UG49HvbjziaZU+hZpZQsZBHW0dr4tacVrJwPrbDXjRPWyy9X2iyYngI4r8oRetUr8OgTazZv
2PGdulTDDrdfb74DDFAXtjesMsZHXXzzaHPX0QSAURpuBAUbmECPyiCHrHMte7Gt6FynTrz4oaEJ
zuWEDNGW1dCur015nj2PrY8UNhOtiLbdox7ER88Kd+1+UqiLUQromqfXEEji4K0GuM2ANLGxPs83
MVHHTf08aJLDK++P+ES8/DB8F3lHyrL/Bh4y9IbjyCpcSbVaLenlz3BYEwdsCAT5aZ/hxN0XyYkW
kL5wNGlGZdKqJNrnX6iLW2YOeiLQMobNC1fUhsHGw0HC10E7l7c6j+fqwHw6BIFJlY6xKcWBmEHB
IkDmZB8+keYuLZvFu0Z7J5hb3khh52dESfcUYZzWbRCxRZoZ0P3DomO9lEB8jGINxmVhDPOnsrdm
axPfCdl2Iv6HO15+noIFe4cYKKwJ+ecaH2Y1Zs4Xztz3/Ekw4SZd+srVQG8SO+rDBFvGMsuCO2eW
ydMeOV0Iyhw/rvHP5gulSJYhVwZ+WijLnQ99UgvsFbhRXneunQMDb533NIEkIeidP4k78HeyliOS
9CrolCbDiu6X6tnPAYwlmQWBQ/ih8e+sWYIVYK2wE6ne0nq3IL+6KSHtvcFPhbKsUJuolfT5NiOK
nhrMj8ANwkpLXxKp8UJLvj2TQq3EXNjZkKhexlVvnk6No8Qk6trMTs39FJ5Vy1aCHYnpSMM8gZ2z
Iqbbinzo8WqVuXFHSgG2iCk+f1oICdRk3Y4WH0rg0KyiMbNK12kU7vW4DTDl9JVB2VHOUZGYZ0xy
yQDERMZMc4ioy+/IJY96KYYLIIBnS/lX230Lcsc09mQOq1/CvjvHsOMyeerDv6G7DveY4D8JdxO3
Y5rW0bQpLrd6/kRbjAH10lXjTzl00EfwvCrf35u7u+DfpCnLRGaa98Su4Jneo5HatapU3WoRF8Po
kc3rYCdztC+Oo6Xq+Yflox/N/oQwH60YWGxyhuxdQPm5gufop965qVjIeQ1C5yrqmtC0RR7aorDn
Y912Qy69p4k8dREihjPwQF7oukIj9wIQttm0DzoP6XcQwt1PEIhbPsH28gfG4OI6PIm0ZIYSnK/b
yrUxsNbk+itAnBjTeCSxUHitgirYbZD/nH0Ve5EFNi1jsaLbQHpd9RCVjFbaFrkgX6aadQ7SfReh
OhN7fe8F4y8tvKFy8jwTt/AYB9KXrJ/dfARpw4sRS9IK9x9YUhNv/nYT0YkgNmV0WSZuGojMIhDV
xISiX8kdF2PhagUANgS7JBGYw4/mMqMGc+mmHqiWdO4Lgy09AT4KeMC54PkweginCYl6pMH9016v
8+tB+psSGqEdFC/vgxZtrUMnAIfs6KtvBDmG4O0rntE0tpC4LqvLGeS8sqUWvZVnMmEvY4+HtEFO
+WYD9R6IiI9Cf2B4MWKvmXqCnD4p+NgEpCxMnR085rsj1/v+0PSzYSPv9K08hrmydpXkyEJgYic8
3xVWilRqJb6EmwC70oyliKvYJUfaOrR2GE6xr+CjZ2nFweX4Pg5XFK0GpynzvbudAsc+w29II2Eg
w16ipsHFVm8pUoBfeqQrekHOrlM7MCdUAxnmj5ga/nYBchJ0RE3pF/AFwv15XT8eN0qm+oaUTiKN
yVLhGAGDFf6QFV2XovAnk7HnaGna5e6r9hokmFdDnA1lSZHJCYn90JAz5LrE2BLKPA8UYKydD3Sg
5csqMoG1WsZhjaotB21t2NhB2LWqof47t7SIMhh/TjW8q/zpAzPpiUQJLFojuScE5OQF6M5YLlTu
yeQ9b1vI10rcV/GdkHCljgAX4PGKWVEzsIhrAUHV1bj8XsmlrFUK3sg/HauNaAVQa+NQpS5HV/i1
HcLu+0GJhi49PwdzUVDB5G+zmdPytwjSqZolF4svF/zlA2SftaijSTFMXhbXvzpl3xoruhpzLetS
loiRab4xJ+VGIGHkOyghJsYGfiJIXa9AEfoPCzeQEJ8GPlHDLFyZ41y00Ja6XWOi7ktNM3hR5Hd8
pvVzlGE8UYhEYyH1noPV8FhMHAuQarElaI6mcD4jRApTxgDbR4D/G1VNM9D7FT2ko8RXKARFan7a
DttTPd2tEnL/ZW1k1ud8N3PhHnvIOD3pR2PRMAXb+eaVVG8A9Rx3dgitO0OrqD7K7KoatsFR8Ytu
BMbD4s3NdFllDI0IKe1O028LXcuioZ10OqDtfuZok/zArgWw+hcMXkYA4WzOtmxDn8+FtSA/0cmG
sQ16o1JQ9H6FhJJiPL0VJOvhUSgyqrUe5zY5SWkweCkU9tJA3Xx9a0uggwAYzH1H3M2our771rTc
8fU2kIw32R03duG4huz2H6bzaQFrsxncT1ZBKS1SZkx//pn50i6odD54ybX7CzyfeV3pbmpbciFP
lgl62UXkKy03SWl4o7xgn/bXXBcxSZLECQkWEpe5wyBdzpmpSBz4+rYF9GnX9JCvQYo6qyz4tRZu
cP66rcGxS3uRJ4+AaHrS1JKVnF7noOVc2XP7LgwvUYrfZ9/wVm8XG8xziPH+rULevrfv7CL1x2bA
ccD2zLfTOijo6xaFWT05b1YWjk0RJiv4LB8WxJ3Bu+lJ2YxIHieFRNzbZsitvYrmUlAGXs9RjOs9
FkFD12s8i5sKQRNmdQYHTNpO/yMP2XqJdmqWSqc94Egtmq8f9jyg1cuV5gpeGYGOaxXmmFJ5Tgh8
wEVwIyDGXdKmnk2Ve5UcsCSUX2Ju2VZbAmiS8qjgLBXVRLr2Au9sVWkeUyMfRmmppBZbVCiHVnM6
9/VGhVZodKw4JLkdHfLRT52iLzsRI/3b0AAwQ4g3ynW4zf+WwOoO0xudYxYk5WRIJ916OKuTB+64
Ql0FdP9UHPUclWCoXKwuUm9Wc3uRaRawguPSxCka5oQ3A56y4awCXNegCxaEQcGCa54uEUI3GcH8
x3QxiGS2sS41YQeAZk2GSSie5TcWVFtdkO6JG9sfM8aLwfl9Pb2X3mJdBOIJdVG4+Rob4haud6kO
ICIy6+zRWslpzdGb/lbbP+br8mFlqlp1BJgKy3/f0lt/ByfDr1CBJOd9LsAogITAuYataW1Mx2kE
jLIp3yJ5cRll6Uk+7r5MAaygvqbjUbA49DTq8D/1xI94D695cb24eVgCN0l1uHZik6SSuYkCfbyW
/RCEL5z5zNs8VanHmPkcTCraw8J3BppxO000NJm8J/9/vtKOT2hGfcYCVuL8y5LwT3v0sI6fsz4i
sXmQ+a6zLH17Uu1UXpfQl/kj7ISd1OHGnkmjp+g+XTg066OTz0N8eG2KpkkCeXI45QGHFYi8TK4M
I9DTE3QQmR9OBEkB1UnVOejtcpKGl7sknypu8Y58qKNoBVtruOaPMusCK1jRCeQbelHfiWGfqZbH
ibhLMLIhkAgYJ6izs5CTjnKNd8FHY6z8SJYOQg6v6HLUaTiDlc05hDmDmWt89jV3p0hZnalpEWn7
hbpTnWpUVLePsEkg7Tj2ipjYe6NbPt46Mc30k+idhzGIc52lTK9gK4rhAoY87bFWmIMmTR2OIwKZ
O3wrHvsW9r4RH7KbtKo6/sgmgA4LbJhjcV6KbUWmmaGZ67QSprHc6Jh0magxJeo0dkTn3Q7xRuLP
HTZbBnJgO0mb0IJppA9Z7bj3b+Y8Iy/T6d+GEYy3cY+CM5iT2yboxCknuAhxJn4c8onhQCMEAdAR
m9J4wACWi/uwQZnp7At3ocMRoOdc40AvoL7AhB6iO1dlZsqb6NVVBozpHvX53ObII2QvDAiVezGx
G4I3FKjoAVAQeUlwaXQVSM65aO2vE1SOFoBxfoyGM+DR+in3LlzVMuAKGTomHYwrJHqqoS+HRr/Z
zbmM6oF8wiXm6NWj/sWwC+Y/tL+GCCPRsPBfm1/B2wxtPtkUeASz6Lh9VPX3lREegC0KRlvsG5F7
Tw6tlf7U7yD/ykQU5oMAEzG9VAgMP+M0oONRbGzJjVQKu4ef93xU3FlOHqkdjFPlsD7APsd3qjFU
cK/IJc+0WDS/NPjhSiI3vNlZIM3XuJ6fhWJlS4cNb+ZIlE0R2gc4PPMCwZu5aPA2nB25DUYtpJ+n
r3V+g68UECdLuv8VzePj2A2NdcSFC70jhcy9gWHnAXZ2ztRRLdfmmuGcMP+kxMZUy/rvugA97dlz
z9geV9MPw8VWbCGrSlWgukm9x9CPTVXJiBQa1KhyFakxdsItfqsoN2DhFEp90Ts0B94iIL6gK6L6
vhruvs22xyNPkaH9+BvyADkJEEedr7oC+gLoyOHHn8PwBHGXwFl97Yzjr36JkFMo+GJEinchrbaT
S3tlKsJ33ziKxqxRbyhK5wRY9HDzPNlB3+nZn3ZNsDVa+W+8T3lKwGBc1kSsL7zP/jbJQVhKOrIe
Pa9m+QZuBceeX65QfWCGRrhq/xvCVgIZ4duk0NXIeRaEotiEemOMy4GdyOH3pIh6/fl0BeEGQarb
eMY+gouoq+lsGh2NoSI3RQ4cAA0kad/2Fd/IgJu8vMIyumhYURR6D4lO/Lj22ZozbZG90O5q4mbX
UyLlatb4EN1gflGIFrpGb8kT97xbzkhaALDjMDsSILEcCGLrjsbZ6Mu6LPwq+BJbhRxWzn3/H2TT
B4mawqV5rKo5ZEOifw1osObPVLYZrz/BszZwhoJOyALC1mUH7jKSzN9Bebt5oBVcDZ9MPiHbzXIi
cYtZKdlvNx58520lGTxl59P9ypARbPgXO2TxkrKEFeFsSKEWaklGEhiVquT+cxrPUr7E7MiC+gPS
n0cCOk49wlEEf66YWa05OKM/wCcss4HnDrMD4zbusVKoEuUhQL3c7swdQMXU49eUmVVFjkn89TiJ
QEfA3fWDn3FnggMHeNqeMIxWToog7DspgVRGPqac1bFugB19RUK1vIHM1yfXSu1kL45K0x6jHU5i
huPckaF5kFXDrB/joVNauY1N+SMo/dwAStKds2lXJXMeNoNW0WWuX5yE23TDoau1XbF1AzK+edBy
FbTJS9isqga3t7teLd2vACsZYK/U+dtJtlXf9TASvyElU2PX92eohnJySVVV551mCt/R2LtfXisA
WBLpwLLljBQor5VIf3Ouyj9zlGO5uikBWmAIvcT8ClrKfMPAPsNvpLCIHKldkNAc8a7iyDRU1U6o
RkLD9dLwbiTqDh0YPiQkrshOupxH4aOLjTN0hmDT1jNGA89xGtowgp3waLOXY5qpmf4mYY6SSrGt
nrux1rQLWRTlCdne7nlveShGP2nIXnkkKSv3AKlJQL/JNZ1o7f+FIXqnyuvLlW0KVzk7n8X17m4v
8xOI8+hc59cpiYOVSPja605529QWeVir87piv8KfJ0QSD7/Q4dvJzBGBPvcBIPe2uKt3wPQ/xZx0
NS/kEW6tbNZBgyRzBA6widrA52j11c+mfVcjas6CNCnevuoZf6/bxX0ogIPZy+SX1tci/B8EMMt2
reICJgOAEpSMTRJ9qZHgCdggfQ8/rZIwc8JfplfCqXphXX+t5pblllQR4/5dWdaV1SMbH4pLXQAu
TpzGotEyxhnECj6QN2m3WEnStsjPGJTK79V+l34llYs/GV7SMCTZlYE4vS7usO15oY15T8DilbqR
8rxHf2FK51yaynLpQrMimIFdHd1McszRvl1npO9dSQRhVUxAIysRdxTR0kLF0mTGKOG2Gelxq/bJ
9APFAHfTJDisQSkbM4WDQiojmcmwZEogkV/fHgIEtvQ0VOeQBQzuISaFM9CoBE7AET8gsfOHdjzr
/Wt4JJ2QzWQkjrWFgflTvJevP1DNe5A/cyPVFrvcLIQfs+qbJJQQY+7s5PkKBNaWWFYVAaZXmUOr
2mMIcas07PpnNz01VanJk5T81tShHGhPMsbcgjuq7in4ZK2dz644/puRd85ElVAyUItlreVGfMKp
BQBElU/1kvzab+92QvppXP6OFeVyVRySJwBLHRWmFs7mPv5ZRJmfel/1u9igyhthlaUtlq/nLB5a
oUN2IHRJFVG3hgqoUPktSqUKKFYq/To2ejx3HJUTiFDgwevQtAlN+jIjq9zUXII0WTbH9UA9D5CD
FgFVRZcKnB6JiEGNdOjMwKEfZXMsbb6g3sOULtEYSMRrsaKgJ9lAzAsQ4EkLgtg5nyqmSRc9i6S5
Hv0fpr1TkMVmy8eFQ3SnyJpun8PreqX7Px899vpj5+M+FlH2nfJu66j5i4YmhhM6x96JI0vcZDrg
0bJHcf/vWWV7U7YOLXNoo3Bt7OPAYFVLzTP0/rsSqOvrbUIJgEUOSu2MfcJeTIvdp4ujJyicLOBw
tKX1ulA4L4+cBGc/e+Po0BtsLPNt2TFOMb65CiVPha/fGA4HToFzCA/mIoSYEI6WXKSIMlLOYTLk
gT+u6sHEVy8k5hauTA+a9ljN3yQ9crUajZi9mSFlKPtJAeotQ39TZ618VQoA3PYzG45KCXgyBx69
hQUiOagczAVjF6iUDYkfwYbph1JblF1Q9Umr2olNZMUMZTDBldp0KCgn3xZ7z7g1IOoiSsSnQI4E
2fpxoHsBOqbaQXpKnWfTNcTGpqX8w1pThkLqdrmr/czeVbeVzIYwIyq9IWYDairPMK3W/f+RPMu9
n+lJr3wANasBkIslaHKN6REJtudBj0YKSyloTedkoAUvMtFdjTqkADiYV6Qkw+AnK7KQ2GVOK4UH
k5NVKOYta6e0UChSB+GaCOWLrzqomNZqmL1l2mkIuTPIbA3aOi9yveW2aylT2FmfirGBUFwyU7lo
5sePp9ryYhL8sK7AtfunMb6n5cbeepkGg6k9IGzAFpEZyVjsdgo53PNXmkGFtApRsqOPZPBGiW0I
QTxiVmuRHKMAzwS5VkrTjFZYMTQIllw94Cw4Y3dJeNTro/kDEgz6jLpGqSDm+LMIJEkTqDfAjC3H
1PuQ4Gb5LO6pr4Mii4+Ts8vMXEqRIMbNEIwrrjX+ucqNLIU3ZoI0VZ6C6ViVfSsnD7jOz/nk7pKA
B7GgFBc/S2KYCtFdlC78mpEY6d/ewRk3uXaJrx8Gcod6zfWNYtnk+F/rVEXVy7mORmw1an03o2wu
Occ2+jtzfFbHiYOTfb9/9uBqlrS1iD5zNZX/jAmrv3O+tx3n5taPKHEAFBkcNRxqURjtihejqSSc
Vrii7PE5cL7UNN+TqFWaStrlRvLUDNwFCslKAZwha01oXoqOHhcsS+FjPaqOinV/CvN+dI4V2JuU
Mf0ihUlHEUSC1icbS7aKUIfwA7JhzPK3EPjTk2gzqIrsCcgaAloD8HZlIyqmefDHEtrSbZPUurKw
DBjoOz727NCL3qnzWXFD4K+7X4+N4ShJR+ZqsG9v2w6tEa9i+ivA2lefw4ccqLJMKxZP5OxL9PIU
upzPnvzNZ8eUsLA8x24q+70rAkooJnj0Lq1O5qle4QX1OcjqUNjjzmF8Q0x9WywPsQKGY2Vn2ffK
hQTDOrvzrjTfzof/fwdNFzD+D63u0A7C5JO6N+tOHpkDyKs39xQOIL872SgZcShM52otXbJAkUUd
tA1xekLFIPknTnvtJ6pAL7d/LEkYDlzrkgvCr6G6649AO0lBuHDLfzdy6SpviWllJCNiqWMzjNvg
5Vp47B267mdMVzHlNxYlo0stB9Ke6C/eB3smHNptEXkk6plSlB/iVB/YU/jn3dHyuv5pk1rnW+Kp
ik4H/hsEeMpm2IxsoNjaFH5i61S0cBd4TdVxd28nR88UDyD9Oi93h5Jg7iWJSqhnq5FQ2wJDmYKd
7ZCjZmf1oKZ9oR0wVyhKoO5ZJmQ9x0QYXS//tOOWp0RJhLndPTpqELPFauWyVpxreIwgY/p5JYKT
Uc6hbqcc1XRAKhQ+nO+0BZyXqDC8hsEKdhOubPHQamuL4wHJFcJpdZp6tJMCElfp3oNKskNCewGn
ePeQm61JUWdV6GK6PXNQWTdwtEJJXYrTI7RJmU0F9o1yIHqUfbhadFX4VQgBRLFkGq7bc707l4vZ
rVmLrje49BlcYZUd36FBEU6a28CIlvogCAww4ADwO8fbBpOkwnczJjX0GXbhTtzm99HJexlCW5VD
kSwDaDQ2iyZ6Yy1Um5rrDlzgkQjP8rap5CruzPrgL3NmiNGQDEu56uLa7BZL7Qe1lylMUYRcs6uW
+UoOT1kXH+sB3+V9A9S5GLWMHj/0XklsS/4VZfWByU+w6n2rC/oWoCZ6oIocbiwPe0MCSVSE4RuH
WQrfaXX2fNDr99+2ZwgLQIHyMZmXJjHchADVittQFaHd2dObcXMVCPnVU1I6U1Ut3RaoU97kIIwv
7e8syJ5L2dvw1/JL6+L0jj33KaLgHwBS9JjhMH3JqIJ4I6KsvoAE7orRFgd21JV7MZkecvNaEEho
L9LS9FH3hK1xjL+HljKdDN0rAwZV2fq3htbhnFE2oEiSgVvas5nf736qDoufLul+/IYU2wqhgCc7
qsoGoaapauRwYccxcIbqXGXD9R0ZZxV3K67yWl+DY/eBUF+jQ4T40RYJ04RLi2sBU8s/UIaZLhnN
Jjf/xHR1+5H43UjwoyXntVwPyC6YgD9xEFIh/pN9lkUzudNufWjYGXqEmm7ITKyuq1rlqplWp4wp
pDuMiXMdA2+p90sQe+2dixpd3dy3QTp/LU3ZZo6Qev7zvm/Hp0JfDoRYPp+gRoOyxOF7No6/SG7C
YqkNLqLreucaU8cO+lLRr3SyALvws0/2hacBHECdUUiClILOtgo3GJAT6T5+nJZ2P4yDVihoELaR
yLxAbPysVuFQpZhdNviFK9MyClUyxwLLpdsVasQzLGC+p57PBFmhKSSR4FKfx1hKP7qB3s/ItTwD
vuaX0jok3X4jLpCBbZuV60tN/QaH5MpKsHbrLhUNORlqCTSAsJLbdR41ChZrSLtQPzTYNDRxF4iT
zW6WfTJn+1Xv57LStIDok2wRVmidOIftx9QsYBVQUCcdGkh4WSQaVqwwM+haQuPz2NhI7/S3mvbw
IWb2rgsts0AKQommcBlMxKiF2LoafxPHJp3Gk86Yf1afkEXcD1+KlL8sw4uL8UyBUrILa52WHRB3
xGqxP3Dlr+GeIwH5B29thwheOPcu79UyjXglA1m4LEVtc2EnvgN/vuK5+AhIDE9pVUd765cIQ99P
ejsJQitotmfIE6k44O/VoOkIXOKXYJvw3V+6b3YGELlBqXsDCy89kmj3bb2+UuTcj099iY2V6ekc
IohkPQQbihBUE1MKRMbeX08rDh5tKl6BcnFFbnOegMCi3KJ59KhkqPzE2NWhJMLCd6NpBkLhK+Rb
C4GQpK6TgCVrmY3I6rpvxHf9Sm2TbXDy1R2w68V1/laXm1m9Why5DKGB0XcfbaaObw2ik+uZ1/GZ
aMETdz4Lj/ZjEwprDgGsRv3fB61RXI0yYOiVSAzku6wcxZem+oFyL3OysKZ9+pwW+CG66qCNHO6v
yzPImdIo6JnURGSNN8XItEytVcx7ZN7JY/YtRoFJcwp854jtOga5d49toPJ7sA4cBlE/c6Ff5OPe
1ZdQ5hnv4CzE/DXLwqKit2PnStR6PMVTUZmGnCV9uXhm6gvQtncJ4hgbCXiHUSvzNmJOT3xnoZ9E
xHyCz9PD9B5nh12oRKQc+RIhA/2wOAXxhuo/YzMEilQwGpRuLADY0Tr0Xq9f33L8Bd20/BAER14I
M3UCWJu9ylpqxkjQduVyhF3VzX2G0t/IxFVXuFCHqKYG8SOsMhhXBJqnx0rXG7ZcF1ofWLD+2U0u
papCxxlKP4EhHsSIT/jWAoABBrwhnbTztTx37ETrMEeptcmC0/fm8hJhsEU2XxcfoDGgU/0ktSLI
uYnyZncec1Ppfa7GDodwwFbXzFGhA96wFgGIR2i5YprXsRDxD7ziPpYq9sEYU0dN72yUB1hjTLT7
0JUlq11cChHFnXJy6BrsSiiQRpm1nbFEKa+YiIZStQ1uPXr6LAPrZ6ZgKLRkuaN4NzTCom69u5Yr
T6JQWlCy/48URoLCnPR0Ni8lANKNiZ9p8ho4GZSIPTDi6UrExNcMgSpGYY37a7o5/o2prtMhW0O5
zDY8rD32chhAPevJvvwazbmx05f2JdhnCFDSEz9RWLAsltX6h1eQWtbqP+vylQ9jEhUsfOyHR3Py
BfE/WUFEoPZ66Z8zbr26Qgph+uk5MY3O+3ixb6nE8Nad+uYd2MbG/XEr0xIGCG+tl+aKE/q7C1Rr
gpZDZ1T0BMDkA7vHvU+1ppbAz4R5hkb/xOrAGDsVZkKl+krPSTn9vJ9B/cI9d6KCkz2J0d3q3zbx
Nujhwc8g7WnWUQvqr6CMaLUsQjIUDw2SezOqUOhRxDKevfc9udVDW/pB92lYJz4HL60tdYM9TH1u
x2fSfYjnzJ4TKZitNIIdNwG3+0hajqM7PhNcdG3mMW6w8ILEOFVoUeq+MrFGqa3D4w0+NyezgspD
okNn9738SdS3USMBxP4xEl7XcTDA0O/LHDRl+VA8jzWjX0r9r1Fgv63ZJIel2jpWSaLuS7UcfzZP
Fp+1y5Fq9rXqadlIA/CEWcut8Ib05VqbGV392jZ1UwrllUkzaPhmD3J4ww8PlEa5I9ctScjZIJQG
6cRaqbt/rPpVP7dsm0I1TXZ3D5cvKhD/cXj4plhzZJpiyNvsCOq6u+OdETkNtj/VS5+VFyNz9DKr
27qxSRcfEOqGNJFEoiCu1V4/SUo6Tz0TYdon7amg2CGz8vi6JgwP29DWPH6d92Zu+13ubBn+KOID
A6GOtKV7wJoichxiKwceYDOJB+9hLXBMhjzflSy1y7iuprOQKWssSEyDA7YjZt5gJJOJdNEPCxnt
C0zd4srLWGQLOAKvrcT21B0U8ymygQ6AZacNROpHZrD0DprB4TetQk8VPHKL3I9fXhkWtvWtFHkI
TY0TJSweQVtUuLARhLAIvUCFvYUZwWTH8KhBBrFKX9ARFYyPUam1sYE8m9B4leLzpFc7JJCwYz5q
A2BOIAjjogUNrmdAAVXzsXdp8sypVJT/F/e/YEN9Y5ApcFK2Bpgf4Mldb4ie6g5Z2pth/F5yiwjP
VMWMViLMJl0NpUB4mPa43zMl7naAXnp3kbtVXoq35EyYUfY0absLrP9b4SG5yHh2/2GTHkQGvsfK
giKZjNsxLnTIilrFyPGX1nl8pam7xFHVwI79qtpdpeL5XuU6AXX+ny/IFoi+5awJx9aLb52Qk5rK
4nr0XXdNEwScoj+uYp0a5wMFr+oiJcaULRmzmSKhHfGVSE1C+Ek2RN7WbzF03JEnf57KckdsLFVL
7WSt4mPLyf/WqFBfrqmELoMVgMv0EFBmjpCnQrRu5OxpQE5Q2sS/xwQSikzVLQV45mPFI+y86J8q
Nnol/ie8yBLb0YkPqzialZh5hLHCZtKKy4leICtAfopQb43xy6tz8GLEPJim5W5to7oyRsn9JfJO
EG9wnngAgMTDEaepALffws3EFkPBXGnTYN9JuSY7FjV5WZzmzdk8R8Xh2vQxMrgVU0eMuI/YOISn
vxH0jv2n0KGQRPj2o/G/CIZCVclGkOlmVUmejgbcxEP/2UvwWYJ7fJIFIDFGamCjp7F/Byb60ReB
Z0OShPE6EUIZLCE/3Egy693UBjw509EsnAExVnHZesV1yaDqoKkdlWBKzVzZSEZHf70yNOhDVAxB
gtCXI/DotGp2IiwaIvmAYQuRM1Cv1UipnAW6RqfSyMbmWgIJvz3roMATmBQ3BNUGQi1i11Sgbgjo
Dh3gcLcVRVhxtoSsh1pJTQQ8ol2vpYXBGPtzhAN9OUbk62hizZAFoVE3OYswGESZDp0o2Ny8yYWE
ARZv9EEQ2zADCdpIMVuw9jBT66c5DuElKIzbMR4n3dOTP2jXkOjYbcS10QnSwZajTgMpkKt8g3F+
1kpMC/6v2WflAf6Kdnc69Uw4gwmluKmiQHhu5Wz7wkVUnWZGSNIeYyWV8pRFIOY78FWJP6Ea2h7C
ctoWuSO2lJmm+RgIZObsn5JtdH37LLagObgo3dmGCjBCmOqps7Nrt7vaDyvdZs61x0IJ7tsMuhK4
oPugtpOZ4/LWgJEZpBgOx0ehkILyhOuikMbllpnXxprtevexEjCz8zszGd5Uur7zTxm5SGfd+2Q1
nOziRQxhoFX8WHShFEfHUcdmrVtV0PaUNz516F7/HexCoZq9g6ZGoXLL3gtkxSGqQZPTfgvd0E8H
KdycQ96MzeKJ5tX1h6acbQgcmOSpSqxZeY7QApX+lXV9lXaboafGY4nu6Z44gDLoWe0bjpd9448M
f3N8pioEhZoAALum38pwUv9PIFKU81k0kivRHY6VeX/3G7FxPm5AtC5s3iaLegIKFqTPlB1mg7VC
k3t3LWO1r2gaOie+iij+1DwhDhik88364xRSL345VrUGGCqwhjfS273SJKY/xnQSDONUisyE23mq
7ddZZlHsI4VMfE7Frm1TjiKF8rarfaJ1sIQzpwHuA/qmbaX5b5Q7phcG79IiY1LSqVKn/i3/wTzd
PAFN5rvpK8SvXk37siID+qC5ZsnZqkw9BEI4SpnEW/z6yo8puCAlIJSmQzj9TVhul+Xiq9mkWbc8
VmxHoMyfgG7P0sY+H30My9uiJkOnRRciEkLlC9+xyMRGqR/t5UZh9OYTu0FahzPa/GEgu8uNV4/g
cV1aDRiqhyqFf9GFs2sYssVP2Jpzke1m2qW9BkUq7M1D/mdedR+kDj9VNOrYxjYmQaWXKtwp5zND
ye2EP6Be25nsn4TEwjoABuNdf9XgVcT9m2lc2Gc4epc7SXeXR8hE78MbMCt3z6rTiY0ZAAI5LZ3T
aLmfh7iXCFcrI87Np6XTtgUDnw2p/oJ2yY+gAoT8KfOLYYMPb8pADGHbPPTZMN9jLvg0X98xjlbV
K/5agMetA8G5h5y2UJM6x7eDTKyq9tsdcyonPTlroqa/tcFisPOWZ6EPKZe/B4GdQd6ozMcAqS3Y
XCWj2dmrXJZmS2raJTgc0t5YGLn/5980JJw1MzON5pLAGBtUKmLyTQ3bvuLpcGml4hsybHzDNaY/
YmnKJUkT2ZbnHsBnLjU2F30n9cD6TFSDsWgrl2fVOcr6b2BtAm6SLiP1C6Ek9/XYyc0sn9cQ+tDq
+3HhJsOe0/11Om0XTS+nYycGLDDO0Iggm3arH5rZLNFUxx2UrNopEYkpJMsVsIiS5rPpmbJ9Bts5
wlpClZeRIqflbFoEOiE2YLssqVLHzS2AIhYR+r3bJ5muw0t66A+bZKZrHXNUfpv/cTS9yXXtO12O
sB13W7ltujdKP0LfENcvNWSesNT1WlrQ1nxPm3oWWJDaqh3dpmzopmCOLCpACq5ttEH/u6ZCc7mA
DgSBUYTwbRWidfTRtuqefJpJz0Rm7NMZKNpO60fZpGoifB5LI3xflhBFNnM206xuSp7rxb+hzdZz
eM888rTqT7OuG5V/hbuPPAGRZt0ZAw1d7Rt/w1vLgmLRMZDEPmtjHjyJPpWHagmOVWVba9+nD7jZ
m1mV9UBmhahlVhH3isuW61HMoIY1KRR634nvZ5Nw5BQ+t4GbP7NtvwgUndILI22qHI/zWiorGfm1
vWqRDqPBWipuM4g8eGsvKu/qQm3yuy9pldiLDsq52aM6OzqalZJJgaTDy16x90Rust4J4R+hlI+u
0Hx9UK9qELypqByREMazkFmmGaXEETONHl4TCQT6Yh3NCfIHMxxSM2UiNuwjnHdgQ8gdUkXTA6Uk
KbfmEoWwAO834/Je8FizLVtHnq5QHuXPivM/Sn7KZkY5Tu/ZRkXq+w6pninC2C8qr0P5Uxxp2o+9
cJhzT82W1EoGuJrPbYdA3KGNkbjj9RP7mM8VTre7gGNecHPDlmVR5gOsipx4e1+YbDGsdOAf2VOD
mSy5N3XSxCU+rqrKDA6vAd+e7FEix9l8ikOmJz/mZrXUYhcwsXMzq8XV2qsSHsYTjZDXfAnp4IfC
KBiHOGCsMh5BZ4oZvzP7qbC/6W6NMRh52dPS5cQX/3DJTEjOcqKdtSqDttPLZxpkCIOWsuw1XoVk
WXRvgy8n9jFk9Sn89uFeSZFwPVddtzjCm5uo4HIDbgWSOZQFDiOA8NRYoVN7JfMntCvTF2BqN6Jm
1g6iTs9TU+vHPMbtd/VdN9Vk2ebz7NPxtEarVXEdqxTKUSEcQHZTlMB0WzUHPKZaoCXtcMXd8RFY
9xSQYsd+z5k2o33uSlYolOAHT8o/28uyq+pVbEN7dyi2vsQl8nG3vpm7XRoEdwvnNkHN/Qecwe6m
kxyMkiAtyaEy3xUrVJHntJ07z7Vr2rLOiYCP+DR/Q1WaYD6QDTm1f5gMQYUH8C8TmeEnQBIkfazf
gNN8E5kX5XPSA9uRptuo2JlvBLh/li98g6P4vinCNK2qBa3POp8FcxmLBBjh9MXClKjYAjF2rvPb
dlgFkMA0AfHsUF2Fiv6pYZol+LXKCQWQfN7dnZG/gQGTk8ndGOTaPdBxLzmSu/z9Y2sFHHBX/ulT
T6wLcEpS3dxPPR/Ot0TzhqBU3NQJtus98FQPfxg4Th0APDKG87G9BBGtTaxGgllrvmHgpE2hfg8K
1MJ+g4acgrjN6JBKtD2Zju94YqNpVd2JkJMIJ9w9iMcOZJ5Cqrl8EerJTBrAyg76M5ubJ9dZu1ja
Ry8WlIRZ4qUhqPX6oCSfBFKyZO/RPHEs051/hd8Ucu8WECZexYrNqMYehFegxgBwu11oGNJdSY8p
3VhfJ/nhB6snZ8Slj42/MDc3HETs3OcKVcgbJApMHDYT1LhKg439KVuoM21ySp8BXIvYEalxulX2
RY4TiGuqOdFa4urCsKqN/WdmItLwjo4lOtEAJ+CyzS/Qrb1/gF5hnJkKT1+tItNbU2O0lT6HH/OW
bIRGDeDzUXNVsOsxJlbAEcIKH9qTh0WZdZgOVbu7zkX34OwIo/0AwFkGISzasDAG5kN4pVKGiwGq
ttiNLP/MJdJ0fjEUckbrx5EXFpg6vcM9GUBpe9M3I3pAJi/fJ4EdsyxtLZIfZ8w/br/tIZ/iW6QO
sBopYTt4n+g2DOyrhcXrLNlq4bG5tZwWq6L5X6DD9LOFYTZyhf1YU3LZn5e7mEzHuu6enO8U5gzV
zD8y3wnrdhTnqhyDRDMlKC50YTmNX8C3PzYh7U0TngGeh7UqaSgbW92vEe7BJGxewlo57EZm5ttx
CKYmmI2pb5DLKnjLB4UG7OQ1oZiKaXwke3+buhTAKMZMjj0P2CLOaOV9/WH0JT5rRzKPhoS01ndW
E/VtWVxhf43NM0Ffb64sRS67K3dPo60fZF8uVtAhflnfBXLSyk+uNrVLtmTf7S5lEqlTlweeGV1G
YQrR+shSKnDU8s/AAtC9qOoD0NapTqx1n6T9vssD2n1TIuxu2NWLEgEGKk0cbs9+7K29yH8fg9Dh
K97wzjZWXQwjcFmxDAU/5wcYcBbeUZIg5hTd12oDm5sQjCxnGPcXv2VHa5mF14IQWQh7bbdcZnfM
wjqS/bddtGogy6oIVqW0CLFlp414mfV+bYXEw+UKltLPejOaviioGdotVzih3PFvQLva8nuCdku5
nxry6htsCisbkaZ7Tidg0TzxZBkRqNnT/HhjYxQLOsarEKyyhADMK1mSVEjlojFyRWeqMmmwZkgX
B5Mib1ujZL7mXZs5cyfCLz93sNYP+9x0fm/tXWIf2oIdox1vpOI8aONB66gGZo4vxHtWcq9zvmlX
V51Dz54HvSWYo0/wgd25cAz6Tfv+TTX9YeSf2vuE7D1RQUyVs9D3VA0lSt2Vo8fSi0lGoW/AJT8C
wIY45JBolkYEN974XTu+iRURCFr1gxbkvMJWku2VTsNjV+ZavW0VfnD09NfXmu+tuqV7NVPztY6U
lwNJbg7WC1clD1XKtW8cu1B9T06QIdCbHHZnAc4ZT/G5qHXfS6Qek64j1vCRvxaSfGpTFZhGcNMw
9inFivEEC1GLVT46xgPJOxDk7b8nudig2OpiTE9odzrxgNTk4OCxfUrIWMUS3MB45BVXavovOf9i
TYO9RTpAT0SxslKRwdlUPe2mvnkzH1ygCx71ghR+J/AQ65rxgKVgeuSCtxGo1X1sI+WDQwbdPPCK
zhdQ2xNJgGMY62EYAgj0VWgdwKc4CQu7ojS1XcvyNSPRUGMX2ZU5c64L7pZHSQh5UrrV1L6mcpea
RH7leyTEP8PVSS98IzD/QnhOd5QOGbyeQ0Vtk8YiYf73I5O/Hw56tmEk4T8KPaUERXNNov+LJfpK
Wmqehsqf2uykzxf/sUCYY525kGK9cfUmah3amAUX+uXS6UMUzYHrsXhd3UrJf/XBzwewrvGov8c0
3qopQlaepeQDPpfUC03m0nlD6/P1ovvPkxhGGdUEIb3TUXR02tb8onKKWy6gocqhfcKOA/28803C
ES0eUiZr8QoWwOvqCgfnqZwGKXaYesQzW2DZrX0qsSPSGlXCs5e6Nimt6fnKL3yAdAmqwGGmDxer
+Bp0cKNhHJDqmAqW/qPwDJ3j/tBHmuZDViZ2aNYD4e6Q+E3shkRVM0axahjCTxoTmAGTcQXwkpTH
cXaOnaKXuRs1/p7BeBskE7saKKiqLe46qqWiIsZ6OOfAAhg4o5gTB3DHqxEse61wDS7NaojheYMv
AnRacqfiVHV9hutZBpRGJtUpUF7gPSoGCLOwj7/3QL80fYu/DOdklvP6/IsosKMH53R7f8pxsXCi
pbn+kOADcIxrwisHj3lY5sGvCD7hsDZtiSXYZcybFnBXoxX5b+1vf4fOG7CRH38yJjHwM1olqE1y
1+CstGpnHlHJ9HAspXswVTpz7pqU9GVrmIHABjDrv1C6TTBKluXzi49js3hvNgK4Gcmd+3tOwxg8
UZ9jOh6nhRZahfj8VljC4Hl3SWs0BAhEucmlWn3j1HTLOhmquFxlg/GjwMFi7ycQWNhuXAd02jGF
Yr41O971mXJ2j2WYuQPqDzeQ1TI6oaE6i4xm9E77Fa3aeq2ye6lEG56ozESP+VSKd3dnHKt//1Ms
QvkHlpZRc9T+JN3VWwZjuajD0czNoqnua3ZZDLKJE+39CvSdVbQ+PohK+FQi5OuzjDKHpsScqtd0
wsfnhpL1gv9BXH/HXDcCuX/PBrgoQtZWASmcoup3ITK59VfOABN0LsrzEnAki7qOFIn/c5qr+k2O
tkyjpjQONO7rRXzoubm8Hbr8NCTHz1cKQW/Era87Sb4xAkrsNYRMPcMvHF8jb/05hX7hzrWeGjuL
35q3SQEx4Pbb75Rpl0whtu5vfUSX6mU+HpUkk1FTACgq5qtPXZ0f41ZaorAsmSILTYFr9Le7U0v7
zKOLKbfWG3INUgHxEhPS2JW2j2b/y5dSIa4uESntI3FB13yR8kpjsEVaL3uFntujQQ3npiuKEg7O
ZwFyBYoMLTHBOySNaqy+l2elUqaaxXgsavLPG6eNg9x2+dTsWEp2hbq+JL0g5h16zRMsPapuJHWv
2kzgYAkvKHkOelUvp1Z9ncnZRgINb0NDpLrGox0G8Qiw/jIirBKD8xbhHZMLVttu3Qji56z0vWKr
UcLZRbmETHPMeCvqoaux2IwSqaBpkixDs3k/UHftP1WoGAfH8GPgdKnVUYef19kvq5I5MXlksT0K
+FCEwSWNFcdy6SH9vmEPxW48sCuB7+IQk0a0LJ3n6eKasQ4J/pSdlrPgUnq21w8LznIlKNyokM6k
G17hcuQ9Yxb6uSJCZf7ajReo+PfRBTCVkzY7Ul0x8wGfzLwUMdy00BgcxoYInMy3gPHsSM15Dvy6
gt/uIPy8t1d/zkFf2tFughWWN40783GfVLG4XqwwsS07wRbImgZTITNLOqIqq+BpWYbYxONVBhi5
45FjZblb/t3egHk33G2pq4uCNrOmY0dElOWu1Wq7l8W+U2NQxZa1qR8OsELKtv4rP5KwSCmyV6xg
i+wx1qZ9kz25IEUozL4D0pJiwxyPHWhlNha9FgzB2+kXttjzR3dYO5qi++dFt0iLHvgxps9AUPrt
neARglq3ol2XsWYTj2l4au3qqKX/OIjw4LCt6SP0BICUoEmNane0JVt1tkMXKVK5BGoRmfoPLr6O
rcNooP1tvoMYSl7U/zWJNrsloth8YMVl3szVxCIfskXPVr6fsuDqL8NyvRrNTSwijfWFligFccC9
CO2hgOybVhHlGP4dI58x0WARcjXGEWa/zBRIlPAl2e/BeCCmEiYUh39V29AqkvlGEdZ172LyUw1I
3XNcYfirHxuKmlocRnL9DY1V1fWpuxBm1Q4kmPQCEqghJWb+ygvoTBinsYESXXyehBbFbIASYU7d
JVKBw89ngudMFCyj0pIalGZy5uhyr/nQt0ZtHf3tX1vbjLg2SiKXR0XK5sdLzg3v/DTTVa3brFQG
IGe3RAKWfA6Y2lqY8yeDjkHw+sp7iSf1JjtbwS1NtXqUSntDbdU1PdKg9Pu4VQd/i1cLzli7fxBp
L7F/STPFUHm/BdtdNrLKmHHxmzLFAmeaGs63Scpci+jJT4I7tFKdEpblJ2T4i/ACdrtTu5Fnl/rT
O9k510jr31Rfymx7QXulw9j3A/Fk4Ai6jzk8GvJDqh34MAA9kij1XtMGZXd7WSQr4ne8RjjW7Uh5
PMx+yOheJ4HE8yyfgbT7PDVrGeW3beVrbL+FsvFA++9lBnyYY0tXIbGCPVEGdqjo5VMOWPCqP6J1
J9RN7wtpnXzFoxiKy7EQ1MkOLtcyj1XOFU8ExBIWCmMucAZKj3ywatnUleyyyuWQvzjJayEigDL9
vXzwn8EKApSvXLXUytVUaKvXdqRaq6O54FDRsYQGSutxFWrWH86tyYHOmYBTPOlYaTlqKg2E9alV
cdQU4ZOyWWU5PmbCsBY3C4Dkf4KfUgNrhSv+jx7rIaQjp63by3aylFQXDyMW4up+W3bVrjImqu8f
qWTP+kjJ2Vjjx1nle6e/MmSaymaCU7v+sWG602fVxyWe0qYcNV4yMuN8cg3L8lTQjgp9JNyDqHu9
mGYC+X40cTRzGAllAIFMXSy9gZ/Ju8A1Qoz2uiz+2KcxB6SqNuPQNE2YsbW2jnrYH1tCDbfO5lXf
gyLZS/cEjav6irXsogOJoMVaPkhmIwNJ53ipTJVM9qGUUHjcX4OIlPiuTlCsIiPmffXS5WfMm1P5
QY+68IuSp64T6Qdnxu43lH9Cwsi5pfSk2g6x5OfaqWCCc9y8ECwX1X72vswMWtkuA5tVWRkiv5/a
a06rrHQSQYBu6Zw2Lw6Ldq3oheb64TadrAr3TXesCEEKbwtzRQlKcbE7p4yFSPBZOmy7TF2c+B2D
VD++eQDIW+A1H68YtCMz54JbRr9F5BZg1uXGpPt1T5zg0rY9PQTyWtWLbgDXG1G3J7N+y2llTOS0
/GHkB1kPiwbVHz63VXfssyExodzJuK1qrAUnZzHB/A1shea3IcbIPyiF2Oiz+3Pk/zMSiLuuRGg1
60DQxyQewsnHSNeGgDOp3nOPHd4OTYl2u63Wl3yGrFO+LKkBzbH1/RAPacTWh5/tUeMrgiaLK1+1
yIW1MmZlEXs2Rv1uYUIXiWBUcZ/iLAuvKQkDeFMvFEM1PP2CjneOkot5/61zEvlzWxBlOvLQlbQb
ewlViSqhMsAVcpU2jd16BukCJP8TtEw3F2mfKQiGiZgR3FbI2+e1rTmF/U6Wpymd7t9khtHDZMm3
4fZZhGQnGi94bFxttJDwCTSORjheZp5bMQAyTQLU1xs7hbGQE4CY9vRdmT58Fe/AO/nprtUZBN3T
B9jz4v0lky2BzZIYlPffbKOJ4uVXtl9eSKS+N0vplOX/LPH2sLgrjuGsN0ABI4cpE71jEivUmHNT
AwJltNrENxoG2d21tF4SHjtCbdxzyy1pa32fKTPLKz6I4AQ7QAOxk54sT65IbGyAaZeaSt9telVb
KaHfL3jnPhpODWNkSkqyXvBiWDZ2frTIRsrNnHx/HhVwXYSh8Vlf3h+5XY1DKvU3JoAmY3DrMV8w
gUWaHpAjuOcKzhRf9ilKlWN9siKLF2cR2nGF0DA+yqWUf86IgVF09BGlCMCzzFxMVrF/+Vdpb3ua
nnYYagFrNbC8aWHul2iSfTXL+h13qCZ8PnPBGsgnTdFUqR0Kyl6jbyfI9CujdplznRiDIzBxmsNs
to/8Xle4t7iP58GPjmPOKcyPA3PC2lZkztHxhvfB8sUhrMknrWsMV2UxH0TbwGdyHkhKXTfk+nF5
UFpPTbfgacg0Ot295Uwl4pvMh650bju4m8lB3TaA7fZs3G4KHRHcrREsnHkTn5pixgR/KNQF/kre
zjtyvKf+XbNWMJ8VhsrziB6p5izEmP7DaOKdtj3ZFXKonIDE8j4P0BajJTgZ+r6zpoISmjvjLN1Y
iOJSkF2LRq98Or4bKJ2mhOQ8nil9zqxe8m6DxgP7uOA5OzBqJn+uqTYj3NdMRyDcV4gMHYUFqAo+
yp4B9lkLjBKtFTNDHz86tbNRtpW6Lp2MvRpGU0YVm+uWy2FLpNeejMgj7MGiYuaQ5FnDZPBQWcYq
nKkBYTATOVnh+JcykpZiwwbZxDu3EiGjHJgH+YHuonvf+tJ/4cR/b2vJfLOe6ndvFXEXp1n/LwS3
bWnCnjlL2W7C2vEPIM0uJP1tXrYsbnuSksYYQz8Rfkc9vNzsAAiQ3q7+7jklVdhwgozVORK0Y/HQ
5cLf8flu7aLYpPicOjysCByufYh6t3RWV9rSdP6ogx6NbtOCcchbaVmc/znG1/dkwHhAbSRBlPP1
IutiurV4ywDIBrpwKq8KCM43P27vfsm+/vXa+xqPnFMv6GHRpsxMYHLLW4bnklh/dd0ratgtmwTa
KTZFu6c7wv/VBL0Ne24HtPZP7OdfOxBGE6AYh1iBAEirYSs6e9PEXWluwuwM1SNPyQoGqAtJpeec
kIPu+d4ynA9T1fiZFAY44V6vTXjEEMqqePZJ8EnrnwOsNWoCk8QQhqRiW+yMZkx3pwbcNzxVMmuI
TXNzOw7esnE2vlPSCHKY/UzkmA3rCN9315oLVowbUUOb3SUI1P/xPkjvLFH6gBVBW5LFCqoiqPA0
Zr49cGcdu7xGqi8gqMjY1gr/WMYzlOwT+KNY8F0tewHJIS8rn7fNIq5Nsu1zd1efBTQQbo+6g/jO
n/9d3fKXNbHs6nP+VLdGs7z8v7CHrOPh3wLpprPxcYCbUdMsFRpbfg6ZoncmiNhLHvOTKescZ2uL
xP/Q1DLNWn8SnzP2mZZu6l3dYwOd4BnZDv30kLkrCe+uezUovbQMS9/m/GUVOhYupsWow6OWOUWk
Fqt/8a57uVrqyBX3PYx9l0sUo43gNoa5OTLA29/7DIi6oJsMtwBzhBnfovxhLWGX9sSK5lOzjM4R
XHqBA5Nbp1uurknMIO/uZJUXTDDhXxIw4VSzIbQ0DNBOVhloHO3Z4a+i40lxjBJJniJUsB+HHZnz
f+j5Yzlf7qvnfHwFGgZPIjnacqjtKq6QiGkMPUQvobtv6BljlBrhsnhnYYl+wTuwEWAlHTqwTMF3
39kPWeUX2yZtZX+gcuG+fIqCu8HcXmfIAXIAO/inVehUwQvxx0KZUFmVxWObndJ8O6ASTiSDy5RE
S4Qx+MrVkbTF+V+SbL+y77sQiVAdP5yEd3451UEgVdNP1qr67quUv5Hgrfz+XWN+Dcx9FX+WDoW1
Hi55b3Yup7IJsgo9aGatO0m/Pt6TPX8GzLrG+5fNb/6e/+/J8mwqDXWCWIJOI3Joc7vN414+yC1v
FK4dLnqYrUGSB5oHjXj/HVHY5bTxGitDh/LoW4+hiE9X/cJ4IzfnU9otf80M3n9Ezhm7Zf3McnoG
epd6Qoo0Yria+VqLlr0hwCnDTYsp8De2HJl5ltQHB7N4eoDb5JcQxI13SSkZCcMIzU9HBhjejTS1
dlF6JCjH8ngfzEyFHYIVRb6IPQlYj7XzQ9sgzSQIIcG4K+jM/S+zQe0c2CxHsGlwT7aUOgu/bwPv
0AGKnO23yr7zgI4SLRMW0bwz6nUbneEOQtPE84aRe4xPLnp4GAivavSCmlpw8Y4LVSqvxK3ThyaX
glnBfugITWlATYmuOTeQUX2F97dB1qZonJ+aZssdbZ4ayQKYRG/mz6Pvlhe8Fo5UiGF5TmTX7/g+
zT3nfLrcOZIVWz77ixCc2APVa0fHTd7qrqwsXX652X/eog62L9OvptKdX3nYV8N/DI18OXgKFEVj
pBIKYFbCyQgNKt0uhSetCF2IghPLbmRGyWtg5w5z6KE9RNax6P1c2KdoYLJgPrHSHv+q/zoIWlO6
R5WaNgdrDoGFULCZ+0QYVbMi5PHrXM12+hREhJIw2gP5CERaxAwuL3vB/C31QmojKasqnMGKnzic
NVkZYpAi616mbGp977l2hjU0N4lHuQsMt1MlZJt/FdSuZFRCcUqAwGGrnPnDBKZgIVvekbZar1uf
aqsQ3L8x/PckmIVgE1/vK+6WqOcEYbPiLu99j0YNIJsH5DysKmeclRh3u7g8I+pyMKZ270gyJNe9
ttG/cNHgY+hbGaFV5f2z3o32AktgUm4Lmro/o2pWMOeQ/3qlwslC7EXobzcO/TZLyqYLxR7NTUi2
kUThUJOsvk45xDWwp94NkBVLuZowICHZXq+0vk4HpQ319ehLCcTAquHIqZ8q4NnlbCnyn5ce/7Fp
Zd30ST37vzSi5ogr+41Vgj9CK7rJ/aXLotCWIXnSm4a8CDpkgsqQWqBicJ9jqhad6xXKl7EvHvKH
69uBmvdAMK4M6My43cpN/YZM12GwGy1b/iX3vDc6a1nADtwuY2bKr3hFlZO49J7fxgj5VeKXzT5n
iCejQD2aXS3MV87KsSLVCZ1wsjcJa92+OThYTNvUXsLpA9335gZrTxjIo9MxPnBB3eyFnj03WG70
jdZY0Rkx24fcnKzPid8UCp0dWYoCDXL8IYTUOpAchN0ObeiiZ8b/5797WS9XRbB7Mysdm0RAS/i6
jrVgLv9dsitHMpXHcm96I7DfhjatlZ8CfTPlnjw9cOLdSnysDGMDfoDopg0FWsYffIFWxy31jEZ5
dh4qhMj+yAq4kaejfea/Z3RCFEQe41TJ/OKe6p5fllSE0dVyr/N9VLulyxO3NmNkXiWrRK1yzN4B
aswq8zB3NXPA686W4t6/fN/L/PLI3tYBTwJsMxuheqpEyzKyg2Rn/jk62oEs0glsDwJyBBjPz/Y5
fHcJ8xaNMo5bG8LlFzbEtv7tSDzPk+IoenQ7dzeu2UHrBUogHdxhWRklCxWAeIlkirnd69UC9KA4
WFDQTpofRVThJiIo5klVYzUL8qO77kkhPk6doV7kIxg5QAbS9lMxQ4BnXuZc/EiDVHfy//aG2L/C
tevseCf09cRlT5TCUU/xk2Vt+xC+eYbAc3b5mCk8Flf7tPLahaYj45jB0FJTRUti7iC2t6i2sR7p
LX44QVId6iU0VyamSKXHkDEJ9FA+ZeQhL+2Bk8e5HBLzS1vFZungQVlQiwiaq5mPiOYasqsh7WuF
mHiRLFoKwWyFRpwUl45XUv9MFjbLb84WWgrGbi8UC+6pOv/a0mzPokk6KxjhQ9D7cEVsI0T8qtar
KrPcD5NDLpagzrIP/ibXsv49zwjds2BKkaxviynZQl1rhHO6nDmv+oie1r6WCWRB79dZOJGwKP9Z
HMHx1siPCBovP440EBfl8ZCf7DQ58rVuNyJzAN5kTqXpxjOjQDQaFV2jBq73uYCM5IJ6H2erVDot
36P9GNyaiTfT4VmzUooOUlH9r14dOvFkTfI2GA5OZnRhUPd9VI/LG5BovtdkQQB2UWx4LE+ZTXH7
PXb1Yezt5tkx9VQ8dyxlsCFRzS1wDMl7ec+0yl9Sy1cP+WyWfgCncoyjD3bqpXRK2okTAHrUPjOS
nQvZ3i7CPmkzXSejf+XNe6p6b81Hlle3+Pw9xOXorkaK/t68IzeMmRe5hQhWqSVG6Y9633EtALrk
kHG/DK9ezNkHoLraZYO6Wfupnu/UUw/4xjV/KN889PZDtX4IrSCRpkkmlOr6PHcMy9YuQVuOZdvf
gUSQxibXc6kkZ3Mm6J2eiuIUSgBvyD6LduTI87XiLD0wMwd9gtz6R7d0A7rbMgcQkHbfcY3WbytY
I2imPDQdv0OLuCqb5YwqGOQlo6DEYkUFFuYkkuGy4uTfOYD+CXBip+9D0gD3tjk95kvnKw9R0xTh
5L0oqD7cKNtJj7GTQhB90/bYPYR7gA68lQspz/KC4iRXkP74trdM+HOI5GdNONK1r0ISqEmSw3hk
OXhwKU1Rhx4PN7UIWHXEcBwMyQtX3ic7fNFTiE6Yf9MgHiIYINWN976EgxEb7Rj2cS+khhMl2Qqb
wvsOJJ5F6K5AWN2xqKFFxrH1uVWcVZSRmGmLNuU2CLXkIMhAUpDyQyl0Z8GyHx2QAV/vlXWEiVJA
NPLL8m5oAPLMRn/UeStqlX6htDIENxKJYJESVcA2coKVJ7lZ76MlbBslJDENp+IRMhs86Lvbt+7z
wcRzwQxg7KwPhbZijb5F6bXgVIcb2xVoXRT0fKBCEUusXxosnHBmhH/Q3fhlqGSziY4ZIceRgsmG
qXu3iX4GuTkQ0oo9y9q8Lc1sbVGGgPpFKkdz9SoNDnk4qQ1ZM2kevoPASFNdLoclg6EKL3WqzEwx
F6pArJSNC/Oc1saazm5M8wS2lWbw7n9+51+A/7C2PXMT2vTD7W5v+I2uYgc5kXJ1qxxLck0OsiAX
wxtkfLKOR8fazw6oAAZopvH2gX9CJs5aBVaiXDHYAwfMJo5g/y/Qk4lRwCTSOTz3m933Iwqu4Wr5
u9MoUXLb9M5srgHronxLWq8ei2RG6lLUzFxb02b/oaEVp0teu/5X7g1k7U5J1knymchpG4+i7tI4
e8pAt3BaiMbfDtVK1LqY8lko1dez7eH5+gcdKTBwgYrm6Ck2h4V0vCY3rPLQc2VcLiOLk7crQ9r2
8QQnYI8nxYstoVsWbYtDgIVnRMU6T8SykfhYYmgKJZkhswWBZfnNy4H76Ri1ZvTbNTofMax6CbrA
/T+AjV+eBsNZ2WAy1/Za0UmgFrQoWf6eNJkln48leXH9NthP1q92K+AIgRBfs83P1LYRzNahzrXM
M/iv4gX9LOnxx3wrz5LKIUajjZu+gxDs8VmMh0i2UIOcm+qCNKtX/4esolz8uE3Pw307cGuMLmhq
iOlZsCv0gPUWUuJwcYU7iy6dr/XqkGFPTs7xrO7WPhXd/FI5NVjj+KJvnfTZJBK3b/qKGBYVQB9o
sgdNgiLwjK9aDr5hYqiP9en4UmZF3aW0wlcv0VdZjIB2gMfBi5pG7BMT3eYKxngar5iUAFNvYTqe
yrx43IHzzRCKN+gg8fNDyxVT+daCLdCzXenc4UohjlZ7vw5z+7+AcnAwhU7ScvmIocwVEED+5Dya
jeGno8aQxCrB3SDO8YxdF4IpUmNok1v09yNI3rbucyJsD0HDLEjwh5owmkr4tOfNfDWVwAbj8f8d
MaT+gJDLZwMbP59ViOJ3eXh2PSy02PaRCtUXBPShgOVjlR+oCtyKrDHsTEqGkOSsXBacvvPlgKXF
rbYjMZC1eXID/KaKdSXZXv23B3Ddy+azM722TpwYiq1qKiqkm/sQVT+EMzJNH74KUDxwcY2rUX88
b6pUPqXKbWgh8S4Mn+vMNJW23UkarP0vTD5vKAze7GUGGqijVpMupYhxeRYioq5c0AFodOmX5YK+
HUt2qNH1L86qHr6DarRlzjKTZR8T2XuVfVcKVX0ERSlfA/mTK0Pe7nHQcTBMYVI2ltlTt9z8Yg1q
FVXT6kmIM/uehz0aKdmW6TBcy9ClLDA29HGo2i4d+bdyMgTo4GOVhczOm32G6DoYRHeTncM0r3NP
WJEMzOvRHPHXBqfH/xa7dlVVTXHkx6z0knvVZa4CmiAymBTGF9aEaEPfVybCn3cHhXuACtkjL3Mg
5wVxYX3nHW5sUHGt6NiGWcnq4UFtY4ArVke+F9GFfHVo6yffAHHUCBHwh4HE0lKbG6lcldZBdCHD
Skp6v3wZXZWoM7uz/Nze5XOpbvSDU+bt7xA+tWVILKNv6zeglcx/RDytJUcjzQE2w6LRLUKETUb3
AGLQynE7IiBShjQygspsQ0mtKo5answYRkMs96AtJrbF5o+M+tXQmTWDKa4NoLMJx5BgDHlO8nXp
P13fAfWHs5DFsDFhOeTO1ZafYe8E3Bxc9MiwDjPCGIwChxfw/M8K0z9GNLkl70tCtm5cQ2jxFF+8
BAWIwvUpZH7hRow7auTFeG9+d7Lw2Yeoi+jVPLF+81rciDUH+LMGW6r22v3ArdFczxc7p7TLkCFO
dyfvynI7Uuv+nW79EM4089VVTklOMbW45lBtvA/R5H3vakFdUIbvtr+cG7ibhfBZiAGtNxZJJxc8
j/Ni2B+gelCF8yn/BFlZpKX4s/ufO88EMnbezGLspzgvocmMh0XjZ1ok3KskcyTlNEXaLg3YMZot
0r6c/3dIQLx6TFWMkMoQWdSB/H3wLIzpRZOu0tBFTIBKg4a7fkNM5g8mOXd7URb+utdDfRcvVM//
WdE/sxDWIpvsMnAkNRKky5PqHJs0Gv+A6dsLP1SQZPUWO9jzzxsTy+j0V0jBLsbtb2bqBmlmUxx9
s5YYdWGQVwXzSyFVmWCCYmyFXCxJ1vHpRwmxbTWlHVKVAm9/o8TW6pwq5ACgQqTGgug0hSZ7Sz0Y
zBdT5EscHkNmV8mEZA25ZWPIbLWfuUjVr1cg2N+YyCImPp+TBxzetIv3Ne87ySSgcJl+zgQyyg8M
bCE1eR5ccu9cNCYRFeD2KInG4LN+ofb6Y5rErH678/BHtWF7hAouz4xBTbbho6Rn7qzjGHExL2fY
d6f+8VNAYRG114XMo+uaOBPHzm4nL0D5BVtR9lhjbWwH0Uzx15W8MO0J91wT6mnLfwsdJ3MoA7AZ
5t0QBbkpYQh/VvbMb4HC4iII9QJ658UmXuf0N48RoYhDVNB7hQkUWAVhqOBY0tUdZ3IQnIcwBwEw
SP7lBZw+hW3Icx5xVtdw/hgyQBZFRmiXPW7UPHpoA/sCFqu/waprK5hADcx2u3Ka43dB5d94AK6v
bBnK957yjm3bBwlavpwh8KvM/n3LijSUvkkMNfP0xEBZJdk01CsvC/7Zl6bWAMhNammtsqBzx0YH
Nq7mwNhRAs2P9AYwyIKynPcQ11ewAp4z4etQDSYP5uoP79L148be+g2w/uXuFjfhc7d11LnuTRbC
TAjXM6g33Vrjio2i4F1kBiFcU5bXT/k1DCyIcUxfZ09dWraBUejtwz2PyZJFdRustb6Uo6tY8FFJ
gCXHC7TPaO7cRiZbDuHV4TgkalKLgR0HJhj2BuE9FJ7cbkT1oQQ1q+vFPIwMCx0fG/lBC+J983RW
EbZPP/vMOVNVcQJ2RlzbH5OPQ2Q26aXjdY1lUTtQwhl1nAhgjDkgK5sJ0aT0Sb0d9o1E6HiaacOx
Zhfp1toGVNWTYSv/vyl0ALURArBA2ZJydFayfE5JJpMiRSYfWuDQJZwm+VMIEO5/jxYG3XRqIm4t
43Zw2koQqqg+UIXn1O8x2RPDNQgUaXgYH3hBjj70o4vTZ+OSZBnE0IzfI/gicL+x5ShtMfkg7/BW
U5oUdBMoNp+PcIMMmVClkvAZLTBpgjFjm/9vfgT0JxxjeJLOxaMI3n2r8J5zKv4YvBmWCnrcl6CL
BcI/Yp0lfjqfQptctzjHfSk+ywH9Ifc/V06FVfx/LzEhVipGhh/D3lRmlCoI8DIIdHFrOSYEWaqq
PCtG10X1fui+VoGmv5/3ccOgVS7WLPZ6eFrdbZta6nnX17JcKmpESr2U8lY0HAE74nk/LKjCMbcJ
40KJ9l7Kb/0p780tEn2//LpL4gpaJ465MmGyOscjUBp81PUxK86eWrQvmi2/bupaA6ucz6sLmaAq
WGBtJq4Wa0LXMB9yUUBXqnucQiA8agLMsK0zPFZVuWEagVfXjm3YrO2QliHcOGQAe/A+Vw6qPGdR
QHxmvtbrVlUyVYE+RNouw63C0WViKKN91DDgKLzgC9PhUY8lGmwQmsYc3/9LRsCYMzNI2O5edgXG
Cdt5/d/JMfNSvfmPnIZ3HA2JxEAix/+8AC9fZIx6AUF2MIbo2FcHn3MVM1doJtdivF7x+weeLZAL
6Yr6WhAImWcOABSNfI8CLbQJ5c5lu+wcYf9hD/vqqAud9nRomvCy6l/lVQSdcGjpuApD/3KdNwSj
NL0uqVpN8KEzqao18K6vV0kjpq8j5c/pUwh0AKSjunLB/SoyZ9kmBBKjgv+N7P5t5k23q3w/Pf53
EiyBmZwMlgFp1MGiN+zaDJlpGc2TolB1rLPi8RGcmxUlglAKv2O6fKEwZkpVmQh+Jxt/jEcI9JbY
Do7Fam8GM3jIxsMmtDKPTCzMLC0PnAZi75jKwkwaq/+TM27rshnVIVRXrmsYW/JhS9dK+/MMe2sJ
20ULLPdfBja73xO/hu0Jb/Oh8FzaT/zYAEmqVg2qiPI9XaDi3KqX8YsQy5hbJJmeTSpAKrs3Ru0b
stCpHu3mQC8WBu5xWfUn9Qk7hSEoWIgZ1Xv7DoHpZb8OH2O80ncnOTOXYhBz0G3M/zqvndUraVY6
XG2/CP+5tOIJxaAmrlDR5wz0IeRuBzlrS2HlPpHAIipyR8hOg5iuzSp933X4r/RhcjQJPiDbiGPy
Ouu3ts5rDugTnhgI3mZzkvnMSArfEscpOSd5mYDl0pHLU0v07j7g06fepeeDYJH24UdGETCzpaO+
QJCCfdTIoRktpex51fPi79hkz4X94YZz0PFmyDVpOXc70T0MIlCAc5mP+XE7f4BEnpU6hFWwMWJ9
O1eaLTGr59Ql07CxGk+MtuVmxInxUGzb3G+GqIQrhcWvTFPM3Uhc8KT0diHRfbog2+uXwRWjSGrO
8lYpqLFaGjrjLcWx6k16AuiLKf9jmC1TuLEOkV02mKCbAyNlt9BOy6wk0jpfg0dgAYPGcuPnXbgA
m+GNSnzoIlxgQAxQklRQM/xNz7t3WJ1gP4a1K7lOSV3PQEjD3YG1oVPtlCfyMeBpJy7ahibzwWru
wsQ+50fI3IDPRHNcdqJ3wwBEFh0KsYbeCBYfk2QKcPLvre9Cb7GolHn4azN+lGqlMyJMyK39vl2d
Itzpdhg+KMD5l3oZQTcOtWCR4zS+31HXhFn1vuHaIyumt5uhgHz0+NaGzUNDcaFZuUlU2i1f8tQq
KALrW6mhKacVwp4oU8w+PoUvETXULum7c7vDZ0MhEvTs3WpQe+QQ5rjcZpM2c9sFhsaCVWDLPhzF
8BlQLldUyIftKZ3ulb4+4mAlpie2j7Zzc5h32cz49xq0aoA4zNbXyQaboWDNqKq+sGDr4HqZCJzC
T+LAAHV1daznSm6lRvajCbTS0c0nY3iga/qQAHPunhNh1KvvuMQEieizXadPh2NaLuo41pPsyO3i
XKTyTihtLyKEBSrm/PmSFKPK6mq1xDCN//oJDyqy+nDEKpktd7F2ZUJpjrNQypdiA1z6ugeq++Zo
EiWqKVL9yEcxUOJNrRSNSD6YL9y9Mr25cDQd2N5lWrIyPuKw3cJk46nIK5IHF7eD5Ti5pQlPrmrx
QbEKpT55xfzTpQ+sANqjxcTL7M2KUsgPrBLpyBmpmGxqVhkZtrhb9dMXHi91tSOqv84NiLzQZcQy
YsLe/FKEz+2ortMIeGdTMCk6s3yFw30H+bgTjuUzXPRQBIfnZfcNcEesHt3CUNtWJAQym5R/NnJ/
RSXxIoAAmxyxvTr8AZ84vnU3E2KpS60BVYXY0yRa2ELzQbc5Epr0rvlQcHYriQlcBdMnuyEe1iyu
ua8jlfGwyLxIa4za1M4Pwm7e0REtfX92Tfy6PU2GmUejyFqupg5M+E+D0tcAI0Z7wKE5DfX/6Rk9
NP97hzc4oB7fZJ/7koVRaVs2a+CILgl9FoFLMkJ2kS9UsqUpHqQFskcIp49dtg+NcN2WGk1aETdu
9D2Bv+1s0yBtfdM6A0WkzCFP0lIDE8xnKeiuP2yIL52AcPgcuzWsZjsk8N72t2fY00f7NBwc1coP
hMwooNgpQjrJYG1v3tJMRSBrxHCjHu99hPW9Budf+nANq5Hyad6wGJGQhU/6o95DmzlAQmaxzThS
G+Orf6/g7NFPT/rXVleTHZcKKHC6KmOjcmiIvrMQPHDDt/cKsAJJ76on301pG36o+O0NS9+GKc68
3gqmYTT1yla/n94R+3QqMHhd7OLBpACtjNH0veiy+izD2YuURwHGUls/yMgiHkksbDyAqSVLYy6n
0M+zDXsEz5BNrhm/v0V4BZ4KKMXB5Y+HHLivVjlSwNkgF5WtGybFpmDsDs6J1PNDLB+2Bl8DizcN
2WpDy83aXOBN+HgVq6mPJCrgwsetbUiWFdy4JGCfb6vKjHW1lXJgH2f40sQY0ilSIwRYxHbfPhXe
nl57M9xssBL5vffT3Ii1RIwygFii2adN0dIV+sqbC4vjmoCBFhOuh+gd4AUV9THXAjyO/eu3CcLv
l01aBVhHWoIcWyNnLLzzjCu+++rnakHeFB86Aqm/gNznHcZJBe4vbyGIjUC2OPH9/13cfgAQ1cEQ
Hblg8w/FbL+1WKldMxiMKy14skM24TAL5FTE0/ppYyr2C7sL8enNLs6dZ9cDmBeKKvPDpy/qxLml
r/Mfj514YvYVq+duvr/nKzPd+5vFXXMGpWh4UtemTgBW5feTM5S/tF5bccIZwxrjA0lZB5oaDu7a
DTED/uiKQAmkX/9y1z53miGVaC1VYmiXFfs2f55NVOZotK3fB5vIgi8U6ZxDQw3+WmPMdyJUjNZb
Ufmm8+EKp3IonQK1rVdnW7GgHxF8bg8vH8xJhsL5h3borFEGpTQMGGlk/9l6Jg+uzfKRl2tu7dti
5p+97HVz/+LAe0nMu8CLUXL9/4da0VU33kNsZn9tQzFBlHKjEYsoykL4cD0uw8cfBOFfmx84NwhN
dq8ThcxLWosEHUeyuP3RiMUXflRxR8nt5+i7FvcHPFEkNq/M8RPlXD5Lpncg3k/2pPOiiC0vgCZS
BFFNR3YSuMfTy6xLsbi+RAAQrFrJGCig5CYIVz7nWJPbQ6ubFkfGI8jC8hL4IRHVF3c/4Ws8ztNH
K5zrgFHmhOufSyh5vefTRuUJUdMpqD54gnloNJqEWKc6HMs4uTNxp9kXb1fp+vGpVJipDGloCfat
V0nNVP/KTy8rncBPxJ6C2QnWsZlEHkvls0/mJwFG9TWv6a3bCyUGo01qFLx8VL/52z+IHAfiyWJd
qMttKm9IejX54gYSEX53kiODNS8KWhZj9CK5KHXRMiqXs3h/o1mWye5hv03P3DvYukt1Zr6QVCQM
85Feq8EYp6a64hz4+4M65VtLLnitUH0h957gudKdfUCLHNj7oTq+vV9u20QQEBRRecZFD5e17Gdh
J3Ou8s3kdWo/RDRvVx3l8OcJm9fGIo59Ga+26oOTtUU5XS/6wGRz0r+s8IF4GYWSZM5RFJke/QZ/
zsuVXeCQvXJkY9arnZBoippEAy9xl882iylIGX1k5CpsandeFaqN12oA5NowsgF1PElqQwkUt8fe
RwqRIJxJzxttjpsNNkYxaRGTJbLbNxrPd8PZBXXVAP1gnG6s3cbfEytqpPVbHQfrp4Ut5KlTWZuu
PPFV6vwmFA2UCXsZ7UEczYLosb6LO1FMnHnZL5aC9DIMRcdhVrjV+viuc6+h6UVaKzozeY7YJCTx
aBMIpQVQfVLOR77+89cRV3jMpj2R1ZTouOCzGcsL2u5O6Mc836tYVgVVSyItgx/ZBEz7GJbe0nU9
038LSP02peNVlxskV4zE6pSvUULAlNG3gnwIL7xSdI0CaUTLMyaPar3LGH+7VTUeX3FJcsrvLnSU
8Pu4Y9lmXve7WywgGbNQqyGszQ8SHYZ1ozdLKSOL0UcUJnSPOCIkY0dURSrWxcEy+mrKe/8HjG6i
1dY8Xh05fbKhRpdtobwmPTnviPj6wsejDnfMkTTpEAeg46js/wr+gP+UHNjwIREuspX6/3Y2wlWo
+m+L5C8P40lVbkOi+lItIs8InRP68UmWkLlotaq6R7N/UmhrBLXZxa4LK+NoDv0qYmf1a5QXkKmI
s84DSfo8rZUNTVtRaihI9ZdPnkn7Q1Qv43PN6/LGoc4v41b2KCspk6dXdLDdw2+rl26SjJnMu8dx
eSoreXMbV7MHQGoCZRgmzOz4lPChkqA8hdGkWioNroNg/xC4cLI8OQxdc0Zsv35gxAI/mH0onSlM
0vX7zcPvcYLicwf9x1ViM5rwM7d0+6WFlMK2bUK0bgsZ+RQmwXgzc5tbKEqk3y5dBYhezydAc0GC
tFO3AtlicJbH9fH45OY0INYfulBNGgdpspuMxRWeIFZhTWTCecynHpY2WnNVEWo8D+2cUU/nl51H
KeI3aqWuTBO0jb1gxB3fXXOUmUNI+rJ1rpYT2I+RqJd7dF6ODBgJ958KzGihrmHFJg5rsuHNx7Zf
S0gBoyk+OX/Bj6UUilu3U+p8hZR+AjWqL2zIfHNiN4Kk3k5BpNtyC/mo5nLiwU06mD2KWdjJWiMF
itQ0bJ/9AEid6jqoNVQdjeF3zKc77c5Bc+QiFMUdtaD/JZ+ALRYGMLT1ebwDW6NMozUT8dreC+x1
dn+a2YSTlQlkMBblZmIwPXAHOL8y07a7kZhgvbFQP42AMc9Q3wSen5fEGHbcPD9pCoSjQuqvYVOl
L8GHZ8TE+LkAoSlowtj6Mg8EckHMVOhWWBkbAPmW8VmtEnQLkYPR6bhKv0hYrD2+6OcK2mnvq27g
YViGxMG5kQvYU2wOPGbBip9uuPi+lRekSWGoFp9cf9TDyzIHmiASbKIDQjxJaNF2Jq5RNe7tPPQJ
T+lnXYfUaVIwfWsf/fvsM1MbWT0766j5AD4rvKghmvYxn7ojzAHvXMqXSy/D5Mod0Yk7D+PEvDTf
oMflGzaE3up8V8vh9tOhKwoM/rToXQcuvsmeOIIRyIfpmvPKvlSVtQRQ1VU7kRkyMm6XU1KGcgTl
TsR+MZEmJD7mxV4B56xxgJDW/mjY6ad99H73tU1mYcEvtj+PT2ebFfLJuG1s5NuehySFs2UA9FGx
I8UjqLbQvEfp0PPFSDit6SPWsOESxhih3nIxEGttLHjn2Nbq+A4nQZO3cwDGQtMOetG+6A5AqIwL
S3wybTg7WXZAhUU9MBabm4TxQO7cCVPbXyuuVGz/vUGRUcgqcxdj9cF7WsuopYHyEZf5MP15+D+/
ygECulJJcgJ7qJwzUv3hIGJfTYNWqT8RUf5rkDd4asrrEZwLduknPRSrC34MxQRPk8YGLw4dSuVO
SsW/2ou9mIEKzdCmlvbNo0++u/5xuuQf2Caq8AaLdW4W5nLQicOAjs8Gz4Ds1lAXJjTPHwHu3xwL
dI3FPu5ZBj85RU2G0QoF3E1w8KnFmoQHnYF03EgPhHlxmBJ+eDj2l54uGrisHuMiH9D+fZ+Mlz9O
UbfCvd7D0CmP5rEVr9RcKnChlx6wbsRxgnEoeke7zr9pHz76st8gD5yaB8Eecoq4VTcEnYNQ5Nsm
HoENxkGZ0JvsSy35zYUzgPBK2GEeQgJ2KXZO6/r5iXdtpjNfwJ5zcry4BBV/B4VJjwRA2wmB8zQw
eyGY1mIhoQKWFl+druZw10H9MiyCC0lXXlIVQqGSA8RzcWjD4Fv2d6PoBWkzknpwyYxnGBBexcvq
juFiTGhtJJXq+nyK6CKezmI6TiioNMfxDzt8Zh06Bk2YxqXvXP4xI2UYwN2NaGYrJb1LVbua002n
+j0KV4HM3BRg4P+ZCOfBL01bCPfi/aflM3DJKofJWXuHychANn33GR9sWyefY23vw75f7EYQSPzr
EzZDzMA/T/SMtkkrtLJ2RCkf6qPW1RzsMgR6zgq4PbV8lliCVZiBh/tEm7LkXJA9vbVO6B9i91eo
C/gHKFuDiAJZMRLOD7EIlfTgzVjRsr5Y4NsRZOXOtKIusbsERxP1LYH1CJP1yPNIwnP7ZgD+VIgN
8mmViAlQp2cS7UI61mH6aNeKbgAmqNOUuT0NLhgE/8Mzj1llgBnCjK4dJ/IRYiH+rRd2WCQKz8AK
QLcOMkBt3AO2niJhMFrhKSf1f7Wnvniz0jgH/nUIlrLaGyanqlFo7nwLa6jJHp6GbwW5GHrkdnql
uXVIz+ik02fQf8hbtF3mzyausLubGgSDS6d5seoJoQQ3BE+4kO1pgDFdl49DZpZdb+DLpuRMw2Rx
0cp08EBbovftTNMm6BLzM2LXkorEkfEMXR5cnUCPPPj6bwuM4n5wnDBbsJ15cX5KEarGMBofEetd
LI3b+pu4djwMQ8snqBI11r3NZSMucCnXgYW1RJeLckdIaQT8/AB/46hXXKvJ6UYtorpBns1WbIhm
nL5Kg1eJ8YM5jr0Ii5WFWqGdTrHWrlA+7QjrEy9L0u96LfeQSJXjbkF6AlI0P++ANyiMnxf/US0l
s2mg6Fd1Dmdh01vKXFq5agEIZJRRrwwA26/4kkXCI66rBRldTO084rO5Cefiw+HyW+oCaSdxiWlB
/BI71fSgChRk32Wm6aNyTjC9aC0EpzfYvqaZeLgodB60FFQXnrksZDhCAPVbyuXd7usoOyHtqvms
yrmxrE2MWmdsnTYUBXBl5noLvpN7QQCzDR2Ua7Wo6Ie4V55Vcr84WaT6/NQNb+SZHeXX5ru07NH0
WCUID4h/3f4BuAf6e4UmbfjCcUdziYyNByJplFpnQxSYpnb+50UNucCmR4dveWVABCFod0H9h0mu
RHcb2TvUIWKIY1OteV4ijZwvOzPRcfXbmNNGeYelBJJnxIffRwONZuBYTu3SvMlEnxo3fDEFt/Sj
eNK8IejLIFa8iUvKgZYyQD2ZMoU8aT8pmvvDAE3LYZ6MVn8BDNmBGXQW/HQsv/dM8p/iSHt2dfNz
P748SbqBMPhWIJNSPMz9+rFqOZddiFGKIy5nZSn5gZskuwxTmuh1xayt2kOVR/Bi07SqpWAuerWl
wWUknpyQGDR0A9Qi+bWn6OA8d5O9mmItx+S6kckRQxPeWfJpXYVOtJdBHd69caHQkIwsup0tSOBu
DJSLV0aro1yVc4MEcHWz22yUwSJMe42ympFuq3rQgbns/wG66StrGGT19lMMo9GqhE6AQV4JASAe
9Zwl/Ia+HV9bKisCRzz4zXamWQH+TXThg3IyLSNEHx8cU11OKZYX/86aAJY6GWKuM8vyBwNJcVsa
8nyAbgipuPDbQ7W8OrnbuoNv30r2EgbT2xzyuFIm3fU25BpQxj+t1comILgX7rGv6F+gOA+UIPgF
yy1rYEEcFggAIs+QiY9QaFIFTbimMMWrXJCO3Ts7aYzsZw76VifdQPm5Q8o/v5WGgT86hRqLa6cX
OJY4g/3RMTMFumntVWjr8zSYaucFCmwdmxmQI7wacrMYaeTbwuPgt93n0e0FEAgJdJUeMcONKfBU
yHFRAIODaM8DoTNe0zJCjmdadKYgzuC4KuS+zTji+gtYxGNUCz4LQmiuRJWh/vcYi6s8b13RN4It
ZbTySSsIUHByBggT2e3J/HiIkqmu1Ej80AGo9VUIA43MPDo4qUUyCqHsbQaBhCnqK19dty6hCfAb
GDoH7ugMFvFwKaYkUtX6czHfckNV9mlivxMWp4VuGcZqYHVr3cWinW4ijwbeD+V9JMW0DtH+D+eP
kYRLmiCVFjp8V0KkDrvYGNSAbZpsaHCAaEpDxPRVbXB2mhT3siiQTzy96wwgxp708YgnZ8K3+A2c
kFmA1v4ySXaDsZ+PnG7ROgS0B/9xVvdX3/pAa0aNx76hCtrZh7B8eg33KzbfIaFezxQYYgTrlSX3
PaOcJ12zqxQ3gnN4kHUzAdtSPivgQezqq5y1aRtJOnoZzaNxMCfIRgdWk/sViuqgHJaGMrx7jNsB
65jalDRqu1yIV2lapZ7+v7iHGKLtJTEUTMyUbnnzsKkEu5pBjW8tC0WoVuG/+bzdLYZISoFx0URS
SG01dHspNlRAdhrg4csrPgN3Drkggky2BsGNhnoGInNL/V1lq334Oloo1DBp04N7JWxQXqKPyQu+
mCqqeNXalSfBGDJnL1ti2MxRI02E2Fys/yTMe0+0iRLntysIJcN3mY6aaVBIIkk/RKn/fbotTUPy
BLd1Vh7omjl9DgSOThI3zlLaug4OlJJDLN2TlUqdhdMg1M2lp+zPU2PPrq5HBgoLS/oqXl9os3fZ
YTmwtvhcE6wGt1zOef1NocdT2ycs5Jh11N5xlCtln1GbjnG7loyzQq/5cgiL8X3zfXcNt6ixFAkQ
U/CLPlugLlHcNaI2luHn/YawrPC8Y+N0SQ10dcPhbuzUNZulPVDQA+nJE5salMYZHbyiic+2F8Gr
BdBTJLH/q7ZDa5SaS2SOvwlKhhjVVXugv1WVESji0MfIA0h2GHPON+kAYavo9hTFXIfHRUTJBEkS
ohnYGZjAAzWc5xThro3JC2KNmQSHSW6E071tYH1Bjl/ZhLwOqunRkF3ctDxYJZkwKKXsGTAkCsHe
G85ClePU5Hh7qsv2UqlC4e9hNpl2MqoQwOu9b9VGXACm84PD2EBg+RaneN3tRTHuPHZ141hQwE1C
vdgDyFdqkAh3uulLpErXIVyfclOZcNw7nFmtvrNU46cB8GurscwboRDUL3pBrukEXVGuswovhFk+
/e83r9g27T/OpdXwBwuwl9zd9Lp+Cgs+Vo574GC4wUAWPYKQSZ4CARgxLXBpI1LV/ydOMlNOVVpw
BgR/XVRlIzICir6JqWId1neoSuYQTB+qeI31Z5uNQQ2J8mMjr0mMsrShenUbatn+X8vyRKvYreVv
hHlYhM2abjEsR3Rcu4YElcqFEJpC1tyt+d+RAOItEbzz0YK4HH3PL9vM+X23fmeTcELM0/0/TdFk
JZ7FCcTyVM0dUuxbdYW+MSwx2qdUh1toTFZOc56w0u+jHXBls8kypw1FyNvNPbGRKJ5LeYyh09P1
rGbPqr40GYKSCUZtGNg2N0p6V9dm1DeT2OA0G5xBgbJqG6aFjZIjHDzJfz9tiCissqEWJMbf/8HY
Uu/x2ALijdtbjVPKvOsCwnywXbYoUisIqOA545OwxeAeFoqO5dIqAmHuMrfdkzw6nXsmVCzxFc8W
VFe1/GF0Ytg7bjSU/n0EJnUbOgShhlSjIGx25XjOGHean4DP8it77kFc1UBD23MuIT5Pzv2io8I3
9kFtKHSUKtnJGA1kgMBOELeE4eWsOaBesu86htl+gBD/ewjRbKL75UpE3NrlzoOXt8rRSXFXA2lL
f1RIJjapiOahmWZc32FiGrKls9hj7UDE40W/RcJx6vV1ghXR+OCMBMXBAwNs9gUpkl02hBO7eP/w
iv/fj9zlK+7Ppjs88yD/tUmiSmOqN0YNgu0gWMGf7eXdniWbPC/ngWUyI5DacsS6Qqzq+vsi5voT
GIJ4psB/pwHUxuHcOheBxY0g4rjILncvo3obh6b1iKxOFEvGQG7fWUmoqtqeXDaK52UnuBHAbRqC
Hfs2SOpLYwIHn0vFjytIYuUBvSt7SfyHgNG9xsQioejE6qjP1Bgu9hFYSQspmUYXxpCDn7XYvmd2
OrtJXknaJRuepjajXt2QgHyhIK5o8/r+Th2p3SVjv7p9B6dBlnxs9JVuNhGhyTJHHz2VkB0AMqUN
3tvTfsxLbgiLYpGkS0w4SsdR5F8HC9iKDGMiJ79Fwehk9f7ScXE2FNbRqseRb9zKm0ZVHL2MaEEO
ZbUeNHp7N3a3Vn8853kYu4OBpdDheMk98xJ0OKdY+Vo1NWNcZLuK54InLWY99zmRD3PlH3KtxcVU
hLUTo39TUZUv0+M04YE6Xv+E7z37rYbmUgCMqFeuIxtV7zujvLfmyPzvIvrIydKNKm03taD8vZ45
7AwqlwMBUGidD4UmdEo0t0M71EIgJlaCPHpxoy7YhqYa7rdR3GLzwzS8jUplQEHUR6MDahsp7cA1
bdJPvlNrHArOc1Uzxi7GtX+EzTgksGl5jptyFkzU6VJjuBmdqRfyinc45pFdYjoK3fcxuOb5JQvU
RDNoTHIwx36qLYo66zpta+GUb0IBuAi0+Pu23pNebzZuIq8cyZ+ot6D0NHUPIlM6bVobJb91DEJt
wwDKH5ISaOfigbLoiOadM7C6VLK5MOrr6KQY9+K97SVSbijiNOnOXIGHkAbAxtwkk54yeZu12fUl
n4BSCnhxmU3cobhDQVfTJXAmoxHiNtISQEpdRdnrpo114ljKsbBsSZSVVruswEC7uS3WGM8wsqtq
BIpruL+Gg9deit1lBgS5cskYO3PnfhM4LRurSwpceThVBSpFqtnWTyLnFv1Tn6gJfpjm4oCJ7Rq2
Grz5NhvqhUpnkl+PEbS4vmkHvK8ieci7NBu4Eerx0V10BcmXujTWcVb6MusWwSziuhW4wEH2NkfK
vNJ7KSf8Qu/rwxdZUOi9FLHxrn+Fy7lfdRotRFhpwGG69NKlpoIycKXVUMTuQpJjQH+FcY/eQ4fM
7L2IHIaBu4u68b116aV7WFgeXHaGQ+HjReUS1ekas0JsrWeMHlWjNJaqXCOyzFNPJWEMeCkB0KkQ
O3w+IJi4shjRrtTjnc2IDrlsaJrEymfRlEi40BHiLpCi7tCkV1+c55FhV3PsWO/SO3gefPXbpPLe
LXspdfw8cptlOGMkM3ZmAYdLn+IJx1T2jjK+h5R4jMHz1hWscC4kfU6wjP07AXVUhpUPl9z8zeng
jJ88FILYq+cP8wx/DT87OJXeBu17KGxLOnZ60Cw3Gvl1nSOeDJ24KfaVKrh7cjUBMQgGxk2S8yPM
RuE+juadxYwCE6Y1of6eustNJxE4BB6uBaFll8HwUa1FM4x7LlELbPDzeLgMxd4Yglr9GDhexQGw
9M2vZwBJncSDVGGbsF8g2R+NKz0uRPGB4yCZeVSp91gS1eJlsEiCT0gclEUwj2eVsvtaJaJfjxKH
8Q//Hx0spBSOgMxDfbj7rfZI0Mdp8yNMU86EtiNUOygNb8euD8o2IU6IRbmOefbruQnIOewaB+xg
oA8eauGN7vgvnYWEcGDEFbMxlr1oBJPChmACoZ6VxKFJmhE2aWF2WrTQez0d+2QU6GbmrWI6N3TG
cRh8Obe91cUH810Vp9HtqontOFPb1OUP43VWnSDRZlwgGALmebjDi6i7R0ZYbu/J2mdBuCaXlGi6
9acjMSl+AhR6oXb9AT4rzptfe5OAUTC9LU962VgO9M7LeDKGI1aWbS7uTL/OzYytwRKa89SZHq8S
FK1hoGEXPisr0yOcood6sQzcLoTqPqdR1rHn3jJBngKtbs6kmNB+y++0RbpkvsAqM6kY1uUzJ8S9
lidR+IHtSwO0cjlorci7x1yI0r+1Qku7wwyjisLtInobIqBazJabOiZa8ocTeNNMroyWlAlHNNBi
dgXYJyvIc37UKoIRW8fCLxZu+CxXD7wer8I4I7az+jaR7ASsO2qZ6fnatGzEgLdyx9ZMIoPC+Nw2
4LR3r5KBC4dxgDXjapcCwZjac/tFQ7K0jFMvQR11LO9Nay+ZTrCh1lXYhPmuZSv7hn69094fPCia
ol8TNAeltboMYy/seayxODNbpOWYxagEM+BXaWlyZsttGONl2tXe4yXCcKcE6gPaMBpK9LhrBXg7
Oz6SeMVLjujwapMYFpHLTCoTsO805Rsj8bod3++i4ZvPe8nKDVoMppab6QEMgpJ/sfs7fC+kmEbG
FBbRlHSaX92CX8vopjnJ0FMg/RpLdoFevaGsL6z3OQrhZ+uwkCH79gOuQAzOQe5PaZFXaAffoVcb
r2DCFbc9kqkK6k2TytaYzR0xXu3mZ4g6+vOhnbpBG2bA3RZlFbWFSf7xJT3ZTJlC0LinMHdd3Gwq
cak/LH0CbfdfwpZZ0uzA8S4u93ZooNlGIh9CSy7j31lvemJas3VYNaNFgLGHM/bfVWiAzxLz/08E
R5G54ihepaA0WyiIKgUJVDmQAONZa14Aw70Mb02Kd9K0Xz+esWI0jwXtR2GmdOlVstiRL3YqHMwV
RjWmppb/pcjZ7AjPGvvcdsvCZZRZ3Bpa8RxkmFK5NZs2XbQUiJmy1A9KOaFdGZKR5HV4DAtO2ucl
xR4oj/mqcaxNbMPzFYIK4sYtq7wOmMlY3fuOwM5XS3v1Fj0+49NDhmg1dkOJpRJlZ7m/Le2TweKf
JW7VGCkat8UDonFgPfhtX/+r8nWlOXFEb91Wo557g1HFFZOgpGLni00jJI3n738fyPcAFuQQMkBi
g8MNGlDdgJ0FOdoA1KPKEI5Ogz7GFCzzm5ZnnGhmnWNr9qEctIvL3AyleBJzashBREcv+oukbPGH
gdcs5rU8+3HPKXTcfcRIqEC/uT5xkXYjpSQG/WBEH8m+HPfk3CHOfoS1vx7/LIugc7IMiMWah+fF
hK2SLDYREjWrXLV70z3IM225eUxO/cPT//qspAOpsrPKp2uro9fA3i+RIzScmpBOqtHzLFp5nf9D
KqZiVORnmxnKAbO0pthORB0+qSrUS8If760Afhi/tdLBW3fojlNkprTpTLNitkskVqCTBI0vkROo
bbT0a6l8Bg+QYEqk8ji+e8EYzLXGy6odegj6y+Qg5GcFFWSs39iMLWhYAO7dWHXrqeIeH33xM+BK
18Pc3wpqAp9MUpUp8Jt5wPsD++dBlT+Ygf+Csjj0Jd6wsslc3mb4fY9PHB/A0wbqTYpg7JIsudmI
EPjr8Cm0iW7qGix3Y4JAYihd5N8TeECz99dbf+LQNJR8d5I+xvuaP86B+z+4Ya3ozX93f1M+FBk/
KoeJAlm6M85KhIR/AJw5+nw8IzFuCKkvDoHgbOVlg7Qb120mq53sCfqesr4KOBka+RphHPgvxbBq
5S5X7z9Mn/OTva+6CPFa0OGeaJnVGkxro+Bd2+5g/q8SeQN0YMv5DpzSqUx5BQgu00+Ut2KqRPyx
qTPoVEd24UMbtmk0bvp5vvoFmHbM4KTOsJt1ririXY32QZy/gr9Lo/RV/fOVESuQf4XH2bjL0fPI
gT3/DNZfKDGjVmfh6w346aJkYkFLZoPJkJkB+aMwRPDqTD3u+ZpegRb5Oql2i3IgrQRESJXWonRX
4almabSxMWIbi8GhXKcbKmyGNhzUANhQIo+OnQhx3EPxj38H0CmRvnawdvyGohUaWQ7FZu8WItQN
PKLuqgFdJOl2/jWkcr1PZt6/33VOb9UcwcGh9Ospt6kAFLAbbKU9HXn2njutP9e8NIhjXmuJzwSv
8360WXUpuuju2SLHmrmmwGOAcfit7lkkhKYenTNW4vwFJTOrOVzbXrBO8FtTCmuxn4MVA8QFWFhd
8VKfHSa0GjEHKlC+uiugYMGSn/L35R/3PNA8tnuymD+b3v3xKVyYKcFzxtTpnLHHYekT/cCFXeZl
0EhGpfMLpRC5C3y/27f9mNRwYWpnJLhaRhHjNV2mhG+azj3K1dWVUj+OfmRMN9HElw8gPjpp0+0+
JnhV//G1KrCmAOr8/QLtLsEob2ARO0AsV3z12mlswkeyReA8wD9DHDhF03Tf/pcmjd5HtBYH3OIw
G00+3w1KnM01lmtrcvElhgCG9VK6zJvIiqNz/AYXxQUHkd4y/8QdpsiaFPlgHwZKO8WzOWaIduoE
bC6T2FJZ8igzEQtULq3QoG2hYQiFSpOJAsnbHvv4cm9I4Sd7EEdZVPYaYJLASD8Sxwe0QU4ENlcw
IsPK+7jQBLBGiFM4LrgVBBIR5RWxyvUfIr6v03DTxMGcK9K8ZnvO9XIQfIDXcDhzNWxycsWlVPtp
S0qsENDrJZaYFxBmev8xeUAfIg0z5zlzwllj0/8eEgCTKZFGggj2A5nAABWSE/jfNQ/jJ3tkNS/j
We+XChhV/5EC9ko1H6ZuhxWsBXK8TjiClguuiNfTLiWecCFoTkmAWoGhKwRKunWxTuxHehZhMFZG
/6ZUur12ikyG4CdHpCyAiQIYcwtr+3k13xapTOsX8rTS5vmNvRqfxbQo7IlQD1qZIeAaCAScvT7J
Hrx2nhnQeFdKrbEvbYJBJdUkhELcYc9q2Fa6dBCb7yrPdjIR9+4I3YsAX4wihTPyLCC6IJsd4gKi
Du8rlB5ihjl010SHqaNgZP8MTu5W/OVI6D5DzJb1Oo0/s5qq2/ygYfGj2TMKoiP4zR60N2rm5DSQ
5WuF7zns64uYpfdANakjYfspWBgAPp6hTPfsUj4xZ1LNb125gMg6RBnOGYAVZf5qUybiG3DfGSCr
pgVa2dhTKczfcEniPZ0jTcJ9qmH91ngSmJRWiO6pmHMFFq4GAMBLMKEcD1nAXT9Ds2VknW+zBMOm
pSed+m1dIH47Sxt++BdQ9Q5lwsB3g8zg2mMMHdieJeTKFBEsT9ciI1rnJAfvNggBY5KZ4k2FsHAt
3w1EiToD4N5lFrPQosfmejPQEF/gA4+DLgaHenjotHG417xkrJplg95ua0x4tra0dQ2DUriXVtP8
0PrEI41PdhJaq+zlqEGGAGJS45RjA11UXXheQ0efnF+1PhEkZFzQH5tJivS9AuPO+DPGDjFwMOO0
tlU89ZSqdGQt+d1W9+muO3Ul7utfWwDkfc4Khj62GRrsKRwsxHMeanGZQwr/7RW/MKk34MUO/OSM
8YNKNAYE3qkCac8VX5vv7+EXRdLbqRhKEKZsnamRSiDvPK9BBTd20QNeP3TlzQYlYRIon6t2tKWh
lpPvF8Fa+UVsiyi21cYsDXBRmiOA862tna3TbPqKtkyFxGzV/HRSnF0zUINRwsgKGriTe432nwi/
VaKgHwS8EsrL/Xcz/reAVMzb7HzFn6yUoblU3E7KAkQeCk3JpNYMfEazNcFnQBA97s0mTP7NfUEp
6atc3Y1z/vcnEVn1DgMtfDytyaB8g/jx9sVpLVegxsWLXTYzqBuXe/8Q8nQ5e6OPJhPy/8TctSeu
I6Tynn/+kVlASBo/Xer4cGGlLKonsf4IE5kla8WPCSw0i20F9SNZdin3XKF5noGM/IM+UaXBgC9Z
5tTMQ3V3V40GJGwoi/cjye6e3r/ibgQRpTfIWpSrNywFOCpvgsu7MYhiwc8AE9sljBnupA3Wgkj2
BW+g2c3eVbIFi/olh67SbRh1ml5qmjoDotv+UucLPM0wgT+AShpvtLqUQycY5jdB1Yom8YGear47
lp/bWtReQxxIvv12zpGbcMa93o9Kpdzx24g2VtbefGxPW9IhkHX/qUQmr79H0veCGPqtyM9AOVht
a+BqHwB+PIrWRGVK37GkYtW+n1dYB3MsJ46Cr4pVXLhP/hv0WsqKFf6AcAlF6zkWARvHGhhlwj26
OxJRZCzk7QXR1m0WLwBMMePGTT+Emwi4uP0DV1R/F5yUyJ+B/dzIHqcUxRGtSTSXIHME//92IaVu
XYtufuGXLiN+AAE93uOBaGkBQO+XZq3U102TINYSecXwNd1H52m7b9rrxAjG9sM/iRWKinaftShK
iep3O/lbZPUlN1zVUo3xYa7VLF08Mz1q//LQbN6Gr6ZjX14w2gc6f5OZeKOqwmCv4PVQqqP0UqOo
aabHsLlw2fxwHOIg4TjX/OBYTW9y6ipaWYeX7wpXjTXOoiOdkEuf8A05bdgo3BKVMzPCn8+8VRnD
Qo6Oe41J3mTOkF+Y8fZQ1poSU98rto8jj74giu8qZKDdJa9b0WZcQ15m0/Wj8qozv129I/cm91Bv
HtttyvAup3f0vy30af7Qx+wtTF9f5HJGGvVaaqNPunxAf7/qq6OaDI/aObV/CNH3Kl7UCzKj7YRT
JvnYdOCwfTfdHyKAX395AwbNPMuA5g/I1xROqy8wrPW0Rve2WVWqrcvrMLJZRcNh44vwwIwN6nTR
knUL5MtXtzIq9w9DI1NNCRsZQoBh1yomdNkGwBrsEo2y8TJ++J0YYJ4bdK7YCnFCaW4aT72Ya0oE
ztxGoEgUm1ssZqTBvLrz1wCSwk1wKZlco4Dodd3PNJ5tgb5sAmYZXlLFgftCrptZwbxfS19vaieZ
A9vOMfW10PAzmZwW4ZlXSRX8LtdwLGa+Xpt126rCRuxSOSwbVB4wmshfFuVLxo1u7a+6BZl6kNOX
oiFisQTR4f1RQESxSV00kkMLK+9PL131uxM1b5PYo0UDXE46axGvz2cImyydfFyqp1pgos/N2sUZ
31/J5lkvyXG1cGwKir8KDKfnS9ckQCHdSv+J01W8WIHwndf2xfi/oiXgURSQiJS3X9+R/jmw5+b5
5HMSC8kBgCr65PBYEXXDoVbvrFDxxloTBUv0cLXQ1V+lNqLyVek8V1XojpAX73y2xlP8wpeP2n0a
1Ft07kjr9+TLaYEy7O3sDN4jOeXy0RRspE28UIShxMEjW8VD8P187//pyXT4hklPDjK5dfkug8e+
b7g70P5zkk0ZaQmv2MtkptQRXWSNtnf8Ti2hspPn5/qWtY4YMZU90Un7r6o2eEJLnW4Bb/IQa8pr
yoa6E/ThPe7dHyKjinLpaw4z8HAyxlEMpomLcTVEenc+RlrfS/zubZyclnViTljq2fv5uFWK/GEj
k5sa6HTOhuEc5Yv7ZX2INk/ac7DUtEmlFtBFhzTdHUL4yBLcNfGC2461qY6F4fQzM8rB8hemY6fB
deSk8WQkRR4Fi0hQwXxAye72MMaB33Vbl8lXA+aCKmQSLcfVE86I3+7OgLP6rnPAZi29oacqxkUo
LLT3Ky0P4yshSY8GZ2sB4cKNntGTKzExHyp4ZG8HM1ab/17i6NxT3R9o4uVC3vHmgx7jRV+lgqcK
NEW6hKLDvp3LtdGteWysozybsFYmeH7YWhIfYx6qeYDop9s4jnLd3SUonFNG4zWh+23ccm+92ZNf
k8R0TGMymGvWSc7whSZeT7gOC2CrjRjVqXYeRBNN4DWeRsrlwAIECLLlB0fGy1ml2Tq1wddOvXNU
HIsfjMIX3Et2bGqVSKoWuxdn7XGO3lZt7dgyvG4ju96NW2kBooEOWIfQO4uap9ZDvRLK0Rfipypr
Qv/WTBD7qTEveGIUBTyNNJfMle25/qWet0LhHk2twmnHNFO7sQ4vspNhDJIpnccKmpcYnGSmESAw
4EzSgL/9Np5xk6JmT6DH1IlOZOFEu/tOipigX+ekL0A8EUCUM1swJAx/DFdbPcMFSutA1XAtal5Z
3f5xN64+bq1M5p9W7PTqK2ZatJRDzzL6V03xGk98uLhdlPIBGraAGed0x+3eAw6SbFgDve3UA5r5
anORF2awICkQ+7NbBHlGed9F+x/g/EuZJPySmCllEFCnF+z3nS748+BxKrGUFY6dcPCf3/sGnoWA
/i8XaFdpMDfnvXFOdPHjRTfHKyZuDWYSMzKVra0up8MACdd97Onj3NW4cPmMaBh9ObkCWoLUGQi7
YK4tIiHz8CnFoajr3CCaKkl3QL55X/BYuXcl86BPHWTgWaPGe9vxkRmLh9CLBnsXibv/zRAFp/gx
AicZ2SONgAtA2ZKfG6DOt7jB1ymr90iA4PzXfmuT1XlXAJMz5gTzE2CM765Ns+jnQH24FjbcEvlf
qkT89ImVeLtFJLV1KUuiLbVKEiQqC/FZ4HOraXqwJSaaA1FnXLMoRWfqTKbKtEW+1PY7aojToPL5
QFy+WVIdcDIWjXBSQS4vkB944tkMcqx39E0xWLdY4qvvxs4tlBMC7mrcte3cIf+vr6KWacIW6FHJ
BKIuMv6e0HPywKE34ExnWCQBUB8XBNG9CDpEnHnqHBYLErePFljRoP9puIy6W2nQea/7Ygl0hxC7
XZ36tt6WcUtxqpqRNCTPCSFdXX0NzCMK1f2SHha5tikzEftirJXAdfJri7o1ESC1BaDF8RUzCxG3
K0FcvK1/p5DRx7Rf2522rX9h2/DBlPRRBTXr0OxnnW6xq3SiIBZrSPZVbB4mbUg3LCGTbBFhWYdS
CIhYzsM25NWe3IHAy5Y2VtqGRlZpiHU4L9k7B16ygxHdilo4DXMSIIQ7Lh5X9LK7YRHJKFTnH2LH
FZDCHW3XbwvzI05PRbT7av/zw3re2H9bbipJF14NDyIhY63VaN1CZ9mGmrtGDfSTHVGfjJdCPXbd
4izl1ESdgJjquA5MOQVDIbPp9bEvV5NJR6ihpDPZp4JO+tWpt3YxuuGxgGBSWxYadTnsgIEwE+cT
wCCZoPNEV3bEEid4dOI4MO5Q1PpORiUh4hehKZ1mrBRD2VVKfZsQo/9+ytr/GZqqNTgEoaNFCQCH
mHyVhYOyHciwqTMqYqFRtF6sA9+J+PGKEmyYbS8kgllDq/UmOZEZB8OWFXHpneXDvyfO1ist/Bzx
c9TMFFYOXnD3ij4W53LUWQn1/zSFC1Tt8uhyEHNQgO4fkwXecykhlUi44U1FP/p45VSF3p21gA6t
yngZnagdcAOGOy6eJVKdJtOd2ZsSXMhq9nA9Z0l6iIJHKsMEWu0HMsDs4fYbbbKzevG82XloreX0
1qLbUv8xzUfs6Ze4NVh+Yl8HOOcYm6zVKgcj5lebuTsxyVoVlhyS8CHc4pyk4S8sh4M5l64V3zpZ
6Qza89407g766S1RobgHlcdgGGdl0hSxTD9frahPUu1CO5pDIiyxDLwawfzfS26v946XkFpDvOQi
TW4TTSBs6flcHY8S882akqeAfEd8wec3o/Og+GqYIqE/BBA/FE/31OgnKgm+byJPLOZppPMgsDsq
xg0M+6A+5nDglLOFxlg8B0gWROeVfnpJfY/Y0XavsjqOWg2d+wtFYkDy2l0rUVwhnxajgxVu7MyC
N9xpuF6/92klwNRCKchjNuAXZUaZoQpp2KLKDtzvKnd4YZp/fZwDPu85gV45ld9FyPfU5QIaRDk9
P/7kNfVqDTjjfEm/bFB09AVazn3eymbYeDQJG15rjjytbq1AQ6ipr8M+p2UzRXzUo/QT8HbpoO2N
Ew9swbje5OwUouos0OjiAZ3qJxzaY/WGICc8A/E7b6/mgbLzm/ilaFcODHNh3MYK8ROC+Hr3Xo7w
6VeILsX5irXkSS4dFEt68K657qo8cA+14WzMLuEiyTF1q6Cwco4DmSA9zamBuuWqJCNT2ClTzW0X
SCvz9wK2UEUzbsl+SJOVBogqU9kw2BrO8bx1UNevc11mXFzgWWl+gA5hPIGBAbvk543cOgrbI0Cd
dU97VrTueQuPcrbeIaXEyCIUkORuQeaukLDMTmw3HCVoQiujV6QfESg4UDmXelMgO4KTIST5Z/Of
DY7FwPou9/WRWugYKMx5NZCY5whlcuNuzUDrFPz6kkzVTDMBGSP9Y+Dp4vDypI0aN0wsfWDsQ1az
/5u34yxRfUwAFyY28GE1MvO5zkurR3BZnG5IwDz/OUfIQhTjENJw/aLmnXa0rs1jBJupDfYf9gdJ
RvlPm27T3mp60cotZ54JgNw+8xXgvZOQ9EAD6evluzhlocHqgqGfI1X918hogJEdxXUUDDjaEfr8
z0nZaEsDgOTDw7/8DKtT2rUPFxifWfNChP+DHO7F4w1H0YjaSIN34zzyXY4Wd2842JtXpGMbGeio
u9QRXk+uRg+gauw1AlJapbHy0z9p+DRfqqIY2/pABQ2uQELyFIOaiW11Hf+MBoRmnOK5ybqzDjuk
KPCg6FcTyWp2snknHR7i5192D+NhHNfQqtpcSHXHxKSraDl5+PfwPa9rnOzT8+aCvfsdpyEW62lk
QrnbtP2/Hmzb6AhyIslMMWZ76tL0ER24ATnuRbegSxZT0QeWbY6GgI+zoKVIeMtbyWS4RRxux0Da
fm0uICtYWZXniROv1PcAqqpemPu0CedH5S1J8yBujziyCVPxP1jf5uvBy4kpq32k8vVPkKiVwxAJ
h45m1ARMmIvtnRXJEKib3AQQphbPU3y66V0QJFsNDBP06A5bMY59mvJ3LjBvuStmtzeq2fuWF+o9
+V/W1l0aS+Ui6vzl2Js/9/aSYQ2Cj+7/VWMitzr0VCDbAv3FfkvwvYNIooLqQEwlCZxaauyaSf76
Z9d/b7yPz9BXMBH0QXoudZjyNHloGJ4JInoK0vuGKlVoAadQKDbLQZJ6gm4ZDFk7LNIkS2/fo60H
IoXEoI4Dpxu5tRwehL+TzsCo2942xwGm4XZI+T1flDYhT4R3qZxrxZvCutoTtPEv1RrPWgrzRkF+
/NqAeM6UywJ2UY0GzHFZbxIkQJ+82ouFdwJ68mIA1IpnQQnfInm7AGRk+GAUYLk5DIW4Be18m6+V
8zRiU8WX9LO7JiR9x3OacIn37z+TuX3jv2oyV8QwF+DY1TSCrhg3lYhdhTUFasKtPDYNiouZWlug
g65eYmFUQMn7Z4UKBHkXtR5qcUN3codtdo7Zps/n23qMwzwmTvVMYxcWD5PlPk61jrj2TDrLg0+L
vBFduDqfQCeAw/+TMP6++Zhq38jQdGCNRD/hc726ROxYEnyolXJOQG/R3B9/niFNSlq3BooLH6xs
fsPm5nahvOaeVg9zx5cNhuZd+TA1otBEb6b4ALN3u8lPjSyEFKxHE2vyGU+b09EY40sdPt/eWkrB
uX/N+gp16hucALsW83pz5Cz3PbE+N43hU4cZxFvSA2m7w49utdMCERu9Dypu0MWnwO7Cx2KSqpNy
BjcQDkgSKEfmsbP/IT9Wssg4f+5pfRSlzxfRD9UZTjXuiGEzHGCSqn0qVnssz16jfNzJFMUXfcrX
mRBLgCRj2IX0Axox1zqCb+LWtf+bGacLEm+WqZqBv3lCOa+wptoIcb4JmU+RnVUppS2FV8Vks+tj
WEIjVKfWCKlY1l46nLx4rp677fZWTcatCEl0+Uul6JCe9qkLDxiorb+w5FZmNG0YlXStSK0TNHh0
8IdTw+W7Qjh8zRxUBv1ijW2xYjhVYIUV9Sbfi88sXOpHufxacs2vgXkiRafNsu4+MQ3MzVAV/IQJ
8cBbdfC5Cjxibao2qOI6qUq38Z62TETQuPQIOmDFZN7sto6WKZ/xzfHGoH6H7+vVS9Y6Uc/ze6LB
5gRzbNtk5SUPyXIr+//alLbTUjnxTgwkbN+mCge3Aff1Oh7f1Xa8y4gn9TucTTdQnw86K9d019KE
kL5uKMsjciZr+p4yQHuV+DN8jmDEo9HSXAFi8oMvw6+FVvcj1G16FFBSTnnWSsRIYf0oFaJT8/VD
JeCtHYu5990lp1GPS000M0fVWoOEOQVVykHRP4ltb647I2+Ri0NvzCH0eq7P7+emLBbe3hJn7890
/8ukcpzBibnQTjhex5alpA6PgHWjxwxsTX07aYANZTcQnTULklyv3lXb8WwCPrLGry6aO8x2FEeu
rTNUTtVvdrlO8WcsLVl3bjaICC4bv1qk/tUrsoODeN05+I4OZttlorqAJwriTMlMVqkdpUE8/K7p
Otc9GU5GpkDyeFi5FVCXKTrSa9IfYX0Va8huAUZib1VvYkCHGVeiySTOxZpi39u98OR5fnCZGc8Z
uMK6SkQxKwZVQfi7kq9C/ShBe6ZPrioTWeNf+eq2anQQ2jbWL7ZSD4xjjG+A7ZVPEseJofkexqbs
BySmJ9BkCCrgWpdamDjvLLDM0htAfkRuyIWL5d6oJ3IGZ5X4BNywNar2iBxAG6FOJjS25D7r3Uub
WiJMYN6xsiHanC/C6+oZ69v5J5eOqvfgrhoB7CZMPAzzBk5HDd59EjxQGwXXdzzsONSzQTyTmaM4
feEyetMvhbwX0KxRW248aW/Zu+fFN1uMSesR1+bJxjlPmREaX0nU/yXCZll/7j+nV1YJ0utkd6pP
69dcj3yTG8NR/OIISeHrctQgvar4npbtiKgEX4JYVVZRaN8ultgx4oBTnIXzxSmbir9/9BNWpJz7
vypb+av6actu7bMBRUwAB5zgt1YozN+mGTBkxlEHgXjoj29Y+5bjvyru2/5UYKVB8f9V2Gfed/rB
do6fGHZTHdV+X4N3j1r9gynKvlBrRfRaJOyARLgxFtSRkb+WKvPk7MRi3hpikS9d8VdMBClInqdH
DPdJFDrG8bdSwMz3D+o7KGAt7d9cd8/Yn1tPx9FyWEk/ia/OjDFuY8hrJrS0Ah+DVeuZhtij8Qrd
8hXcyO2Num+mV3R2KjIqh3cpKuc2Im5CvNtLy1bhV8mKjeX3JlPg7Sfp/hXnABRXk+hv71qQEv/O
2K1QoL8TD8n+YrU95PLgRrVeuCK/fTEDAQLmZawkIjDZIooDI7t5ukSTydKHjBhE1s6kEz1ogyvz
zNnz6fIBQjWHUYEbghQYHWbVtn0yM0JRWwGNEWQcx+FEtQMwVwT9jqjPhtR3sZKO8gxIILLI0iIR
Flzkngb+E4sPnKBLb9bwK7TFWBsFDbLgbniFGvyWypgy7haKdPLhG5YGmy2mCMCH9R+uog1K7yGp
9pEhmddUMHtDsaC25vBikQuJ3FhwGkhmK2OG2h7dCT8ZK8wwqiDr9BWehYZj2xLS3UUB3JW+qJBC
QjYkv0ujTb8VbdEzsvoI4ncW59wF5Gio1H+dcY2XOU8MWhtO4AUxn3wQ+eKx0448yq1jy77sADND
D+TyTDU7XLU2m9keNQJZsrmEgKAM+/RcW13u8kkzJPkHKuRElSIEGD8QUJjqqnfbeEREkejnz05N
3RvbCrJjT20DmL8jzKrzLAf0cmywTb1CkoVJcvaSsZcphx2C/maCEmLHp0OfGZdnfajO5ZqoewkN
hjay+imeQzPgxqhlNhIoza4JtPhhGQ1VhI0CubWgCJhNs1UXCbRSp45fUdrtFhV9ttAsERcyvwP4
AmCDjIq3URC/VAf2wDM3ZtJz77QkvIqChBQs+Pz608vtGCkMyI5EELQ+Vbidlefa7BU9FWTab651
0DZnPxYEOAhzEwakkpJF9NgOyqDyczR0ifUQzWoOpOqH2wdnK3SE0jHqdsyZtPYuUexT4OUMZ+Fj
SHg2F8Gaz6x0EzVGeVxs1j6b2lz6T0PXMG0SIjGrUzbjK3tZxdnj87P+i99Mx17JXZrLGejsUdxK
9nl9Gj8vGzWKkZRCS2oEhyJwMv3Hf3Dt4Zadd04h9/6kcIuEQ4LAU/u8GSVqNt4JtQ0TksSKBlDQ
woOI0tJD7LaV1LD8Mka+Q28XAaRfrjv/1JszxbAb5M5hL7smu+if5dreg4uVWlY/jHX8mlW5UNgB
sBcjnx278LB16mM3NoFCMNQTOi0y+7HD3kZKhchipkGm3xjbOfon19EupL8WnVpqCQ1rEE0MTjBh
1WZDXwjAIYayN7meUCWBL3fj+/avONeJLFw8r0WYWDHrUPpvKxJLpsEzJ55X0Yc9LsdW+LgOCost
y82UwVbsn+88lGHkAv3vBFwtlabII9peTjSfz3Y/z1Mwui8fH6qo/i+f7tc0tCkkgrnx9i84JANH
3GYkJKvMmPhvVT/DSarE/AVo8kxp/MGv5YMfSNrR2VVhhq5xNHYOaJfMxLWXLs7POK9dkGL1pX7z
wDQIIerTkiNNlJu61DFW3Xy3TreghM5BgsozPaxaDbW7XMvpkLwAiYvWvieIwtEQxg21ftHDHnYG
pB8JG+tc1kCJY+4t5fNr4wChkHk9Wa7GDZ2Zi2l+5QeqS86a6QJVF41pCr/Oir1eUSlKGPY/8i2c
5gbKRb6TZrtYaBTSCiwcUJ42uW4JLgFF20qgP+M+TpCQIOrSSy4BbGVp5+UjwyA4ounoVFIe7aGn
qumOB2e4VbeDrnbUKIMOUJ5xitH3yPYh/CKmS0PF/5Hm4MF+17pUxGjQZvQfPSAlky0CY6/lamTX
BWSnlEea8z8tFYjfnd0A1Ms8zLT5cZqaeZjZtMIv8xZIoGKru3eVNUmEGBohieME06DwMlSnzwsO
Oo4snfxs4e/0X+wNZzZKEsU4YxHt3TcIkH5v1t+kvIzCF9SMHh7nR4JhoXDBYkv2HgYXYmO/XiXy
YJpZyA5k+kdNZwRUzLMwu3L62C87HcWy2Gek8yiv54zXrc6dLwy9CCsvl4T3nE0Be7JqrLxUqphG
YtuQS6Pl53Nc4dO7Wcg/KqExMFzfhPpsNAJ+rtnpzVzxV3qOQDQos4robZli/HDHvD8MPs2W0iRQ
FF6wmXE14RQnEwgvF/Kf0SuMcWAAD0Iur/gSmuGRAXr502sem4U7Bb8O4LnzEX9qEeudEv4M68KV
w7jYcSLu9Q2PzFHHUSX+t5Zgbedv+17TbU/pNlfGjU0IAP0UYkWNv6wmIeCXwY+hKUuvHaGjvCwC
N7HjyMpXKRvNhiznSb82vyj5l5Zb7bfC9CZhVwvQSKY1nbCHh/FYmZ+VEIYmzOtd1IHcyRK3Q+1i
/XETE2eyB3iwCfU3p4XljBTksIzsAnfv+GFkbsodNqgKzb3upwlPHoWmRgrLJmsMdDpPiYCpun/M
ZvSTr4VwwU3hMycbgMJdVe+nzYgl660Ol5jJj27wN/WlVifWP/HESORut9WfEl+oNdQgxJlRy4On
O/NEEot00wC+84cNRhSZb4WP89HqNkO/+bs01sc/v3FE3ekBsuQfQSJ8HgPBbZJNqB2MjMktMlIg
6sayk06j5yTTUAhJOhHI36UJ9xlSfEiKCJFWCNBD99ZLFbB1PzdPYlfSqic3US4N4TZ6PvHUCOKS
9noxKREyrb80aPiTTGIw9jDSDoxIbsagqmYd2LcyCtG0vtWIGfQDu7AmoMR+M2yDRfiGvHuExLxQ
s0BTAtLibcL1J727BTTLG604p1HHP0o1i+qb+m3PfWssFvHHt4lR5WUt0G8T8VywTjtv1WhUVSGB
sP2kNbYYXMiFqniGTTkrafQherKeKZEK/xp0WSxfl0UFmdGCIKQjxs9wbWYe5SPMAHO9BY7JRvnE
WXFPpHMSGnL1N9E7dVM/zVHq9ZlqJyALVGJB3LbVw6abVxSWrp+aqu857mDYhq7kDZhWj3tnSdp4
is3RP06dJGQwZtDO42nN5w7ZAaiUqjblTI+533/dBs9QXk/Utlr190KyVGeV2hzFU8/FuOYVH0l2
MCtj+Bo1UTkQ9HdfIq6zfa8vPySeNADgIHkh/F5BkvqYS+N2M3YVpPTga8os4IbfN1T+zBI2mmDb
MTSmETJQjc9p6r0lXgw+yZPWz9fFpbhirzdGIh0FjurYSyxVBhlD9S6XjIPkamfmSSccJrwNTYkM
XlzOSrGSQtI2BDmF0scU4R1sZKcoq/noCTshBYOgGK+dlPwMZ6Q5m1u55HflDk5UVPTiTN2L+pWx
20WiT8cIFVovRqFDyfT/XT00r0yFo1yB2cukGtKiTB1469GBzQSQz610kKLA5n9StjR5EBSGWnDn
5kwsEZOnVxw507qPXds7SMIwld06U4jBbN7QzuU8vDe/XCfVjiGj0ZQPPxmFzZOXtCiylLAdWu80
OJ3tpIMQh8g8B5FFYYazWNyrQXWavTsLeVwIWPeEYV1etk2aX8wiS6zmbBXDhpFxhx8vMstiqXsc
j/8u8vBkGROTvGAWejGf3XodvwIjk/SE95CVCPPhuaM0TPi5auyBDSkdq1VIGqffo/99hTdsEsBB
aTMGiJORBxykZ9/AwBqr0DwK+4IvSrfy9cw9Nh7GycpYUBo6Vj4oG22xCcTAdivlHsD/N8xsnyCs
4T9/ByH19fuOuXpdnAIWMcNE/IwsCPdt6DJhpJzihrPOghAyzZhJ5slgtINRkx6DQmXQruoVJlfS
4aCZsLTpddYwqxw1UK2XtxSwbBS06h/MH+nSKBSR6tUXJH4fa698+bOdxnNf8bxtGLvAdNKvhGq9
rBNUOmv3CqOaKCzZazsWaFeOIUqVqX/sQ9BovEhYaNyaFY7APTJNTm05AEUB10em3VzeT6LNkYAH
k/ypC5nXwGpgjnXCXdOaFngtk1ln3Ur/zMB0X2YPtBDPMZEFyTasweixvfnhdKQ+OwlfqyEb1gcO
UyWgC2qSH+7SZYiT+BkNjS5UWpjsdDArlUU9MnfgcU1qX5mFoBEtDG+/Dd6L5xi0EHToA4PouBF/
XaknzfaL5+rqNG4SxOh2dr0yq/Q9ydVGTp9NGsZm0M/BuZaARCB7du7NnO5/LeFEgZPengXKnDjL
Zk5ta9noTEaw4uL645cAkBMmc4GbrmdE6wRAFPT9cxcNjwEofSm7VCUJrqXFU0YHY+s29icaRYmz
E6qxjuJtggDK+ZWpidamBzSbPRY1ipMhIglxbe1n5WOLUKQehH+hDB82MaA15DXf9maSHwZln/cd
wjKTut6V/yuB3MtjEe6bBXc3RI9u7LdpByF5Uo8mPmqPLhm9xaXCCInr9a4f9Gw+ewVnwiVJomMf
T803xxX5mDNHPOWK3n6YZo0LCB/KSUfue36Hl2hGHC94T+lPxvv9Pz1Epa1aEzXRFAKQHaF15kAu
9g1rugqDgz18blmSJLlPPnQRIILw6JJNg9rAPCbTQdfwjhqaThNVPh6NefZmvUGM42BNrWp77Y5T
YJ2qEiYmhrXy/KRPLQOgkClSaC3JzTpK7abHwnd9JJZcuRCw91/SpuJsYFeXwepxZ/R8JLbiv7Vm
EsH2mGPbukCPLIDrx+IHaZq2Mob3CDPZ18FNOYzHEHiq58H2cqUX+g3VdjxY7dGL5Ff1vdIak92k
meHBKcgriJNAfKWuSh+Tix75wlCzihSEaSQnSS661jseeugEFdA1FbN9Uhw8ckaeTaq2HTvDL12w
mlt5qzZnVBywL0J4PW4SwkM15dcay0Bi4iettLWEdrcP20Q6YAMwOtq0FBotkT1o7eKOaL+okwBq
WUNZAXGAvULuD2GJ46FBf/RQZsXOsjqHgKm4nd+4hMykvOGlV5cXyIaGj3zXwYn0UGTIY0CbW1O1
bRunGgLSP00KsJaZcgopwElPQUf/p5GhvEgTRcU5L/thY4q9UEYLt+MO9/PafJfsWuPy0tP3QnEc
ooIzu2uicEFIeOqQ00HljRKNWctHp/Lh4CmGRFzUfkzQ82/r92M2Eo5ibC3srcFMDugu3HIF0pYY
TeXIfKEImQ/lNUJrKvb5JSNjuAYlYsBHGdOiCjVTOtv5imUhSslzdwjYq6vpYaK3ym55sXc0tTFK
Hdyv+iFt0O4b8J076C4wFy1Ges3R1tq694fTka72oFMrDOa5oClJ/JclV3f10PGE7vPO7hMXlLb/
JVI3xFwMCNsLfCXcmkVpO1WTiuZZftdTMGTizKZZs1EHrYIHSLZBwtETeZ4n8HIQ+tSRAvC9Ptvl
76eJ7PKVshGblhhXeTxVceJgKeRSSe1+XfZs6/CWTVmNZEI7vuJfQI1D35N8pnr5rlBBZ/2NZLzA
xe/1uU1ELZ+2CmFa16AHQAL7IQTg7eNpbj+rdUhscbJQC+Roy+wV9gSYJkF0lv3JufhXW8lKmkoO
pcxFdAuS/rbuRrW/nXPtnxTTVWMXTA40UTPzyriPP+F6yUYuGnUDbWN1Zgs+9YsJuNHL487dgLWl
MSKIRYp6JSusoCQ6o9R1zwrL1168EqcHjsUDKPccvKADm/YOa0R5Nihn5a+AWURAJlDCtmxcdNrc
oiI77SlNS9Ah0F4dkyzl1A5GvMeJkti+XU7bSlZG8krXs4nC5LGIwb1TcSDRSeWGKbwIm+zLqH+6
7y0Op9G6saeQqa+/w8H8o2P/p/0OecMcEwT721akCuhaBEL8cpNBZtaVzG+z8i5znug2cRQDoDmj
3Cng3gp1Do926eB0teznCxcmR5hiXJBr2kVm3ZM1GKQs/RFPtUxVn5A/tGoZjhY2O4CKVURIb6P7
+Db2CWQ7YHoCGz0JMY5KvP0ZbC3Bv4r+mNEQCRxvxHdT1S/KuOnAoQBXnGyFO74MRlHDXj5UTa65
X9tisD73YTuBXG44XMlNdjJDP+siNePO9OTa5yqByn28McmW4SYc6+hnQ6Lixbl1FplZB2HyT+es
ERoMKcJNL+sYATnwDQsDKsNj2YYrs7qNlsRLRgj51Nmxp3DpLb1EivJ+dsPw1Er82/hch3d5KF68
nRIErr1Ki+L6chLAI9WAeP/Ssliz/hM5zq3XAOTe7eR7mIMyia63mwalc4cHU54RGgwfioLU0fZN
OcoUJNlaGl6MTRH832tQqWddCNsCccbAlN62MOYZeX6ABGUrKqYZkFfXfMe4StMw7UKI6jguDLOD
gdhn6ixVZbnt+5tYK0faIsdsvjdnZlpKPjnG74+cRGMtc3KbD2czwE/SMhaL0egmB5Lr9XPZ/KEI
tshMzFJ/9j8OlNzhvEX221YHcbpBsh7pX1ILPxowFIr1OYKsVV+OnCHeBsqC326g16R0LOSvsX71
6mJNBu7BZF9QBXA6/jACoSWlxRqv9e6qJxtzssZyOSCsAXPGE2TGo6sbu4sm06hgUf+quD2O5lz9
3jmzJNAPkgnzx6HHfY03SM4anZei21FiJquNy2REXP/6G0kTz0gb4FO2xmC8gf/ErQcW5GZom+/M
b3OH8kHDx4b7r40cy7LKw3iuNTuDu/Ejc7v6y538MNAwgfVfgjfzMJjq7pBYveX3X3SnCMCY+SgW
U76fj2Z17sjWA+xkNTJOv+wg74VXzILdxV6YmtXwwNEd8cELo+zGP8LP62ZcxukDyUfSNuinr8BT
hAqqDBeLVwTtY68p9ZkA21G4wNoU4tbfXCyOv9tvmLNPNkgP9xUGjVquH+DW0WRMYBo1ztugxi2H
LgiiA1STIRjmVeLyUvxvOjXTVQIfr4qk5+x4jdL3eIOT61RWoqzlkj1IR28fPrRv3Buu6PDYwQrQ
bq1bbwz42WI8C8EdMSDIzHu7HutPTvTToMlECcPYHqK2+DUeicoqrNw+vYbjnDk+8AMcPOB8O79D
/SpGd2578mhQNIKieQWoueM8hK8/kFNajARliQeMGjA2LIC5XVIG7DCCDRpbYYrsKgpkJGRcD8mN
3Zxpfkw+9gRDWaO9Uwzo623KN0YEUkmn6EEp0bPvoCaWKSqGLf75IHo44sx/3nf7PLNEC3bCpLar
j5Pm6YJjntjPqTBqW3x34F6v6Team6bqGVhol6vnl4je7i9UuioLy9//QQKK26TsjFygso5XaAmK
wsE4b8v1za1tXgqBGnIWTYFBc79+jz/lRq+LQNaWLyEpPBSJ8bJechH2Ty2H22YMy+7xNb3Wtubk
7zj0/jfoQDW1eTTVRWsr6Is6u4gTHRPhgkpbcDV2Ve4R2PvfzWDPRmHrI57lfjNURIrBhStSKdVi
pA8QbzdnkXXl5ur6T64YmaPtGccGLYa8McHLUvVcDg5Q9E4bzJS32fQy34QYHnPtaVdsx3pKyNS/
LwznWKpbrwyE/QjyjZxa/mfL0a9zUx8JlooQKAYbXFQfSxoFh2kncQaI6S9hdApF2CY19hZJCyJ6
2KXhv/5vfjSvNCyNMxydVsBK51ID7vQpwtgkaAS8icXHXjSfEF3tjbUYA2f/niCrgKh6uXz101lB
qRlARmBcCvFeNsf11UTuc83zy3BsWDeOyZztDey15g/GM9L8QYRgeD3gupBfcpjb6ATxeErfbhZN
L52eruoo8WGgpR9FcKpyjCBdmFPn4TnjgW0dpk6X3pSNVhU2vFa/8xlb+0bqUGwdy4918lu7ifwF
1R+c1Tk8WFpHFUkEytVM1IxULN6la5bVZ5C29h8ptZgBnyOPjLhfNXT2/Kk5qbcoLBVp1V4h4AMn
aOmCKmLNy2slKWALqdXIa7YLe/cdjymcFIb9CStwkTtwTHcPfyvINBpD46TUSucUPlFTzWPN+6kU
PMeerF36tMhCkI3mb1hE62rZWNweJtyNZaS9UTouzzqD65GDrdnaU0gTxPfop0ghSrST0ZgsqiYX
9pTfJYabU7ZEwryNSCQJYZN0uj2HbozYyzbELn31ANjzNVDXUiYlV04Wbts1Lf53luYIwZOGJCcK
+mvGwch3pExYWSzrNGeKX8RBZPXNRrCE8NbmTRtsIupxLxlSVFsSvWSTIGhX4ONub/P+ZMbNUVuO
5voGaL+1Ps4p02Zvn92CUDbKzcX+cC1TN2MlwjpKeLrLx0dYvEQFb0/7Q44yBTSy/RN7Ablof0EW
efn5gMyQiigiibR/10dqh+LYtZq/Pb97gVNWgmkGepqYjyPT+NZCPjAPFiEcdpCS8xlLH/DMxKi8
TAnA95wsVQ9rglestx2AI5hKbA2SHcaUVEO3bJTdaU+T6YMoXcEl6ug5OEYQwXuPfLA+S1pzW1r6
oF0UIdbpdyULXEHbK/Xco6SPr/llCJwvmAs5NH6oifXTvzC78q7bjBqXjJjDwfCPXi0agsAD8ZAh
K5xqAcJzjJ/QDifpf9M8z1fufRsvmo+Q/05nOp6twljpjm8hPeCVGWcrTspd6olwlg5bYrEq8KFn
1NjDUs7RUfaVombosyxgc5I9k8yDRFxygveBjlUHhXrnDXhGJ9qE3mnO5tv6X4vxe0hDGgr2Va8P
HSPYS2fuqgRM/z+ZDAZ09IRCuxvZYw3QMBi+/a7Rehc7J2t7BeKmQ+ex8/pXrALj5XWNlmuzwc0/
N09pvwsOajEidr7xET31sbwAPAZHaGLwof/vgRpBdBxm1YtvezAoYsSkFt+6eQNvlG246rRBSi3v
fvOfo9K0OrlHU3+7+gaX7Jxpc6wZcSWvsujfp3/XnOzaZLZTXe/2beiewCyqZ9DwUiqDuRPEvC+I
ru1eA2qNtWw2SiHI3vRiO+rEL/yWoc+1Th0C5DhlZzVgvcRNxIdMYPmmju1Rz7AjbeTCZ3GMIN7z
OjkE7OkpBGutjuDPxbCszdzSJnRwmYm5i145riwClQz0rnPNVRDtrohqUNyXN9rdLm6NuXgdgV9h
iE4qDzwy53AaaxN8AZpfslikgGjgJmGBNDJGsN+Qr0jbBSbuMF0PNsg0Y26En8h4URDBfSWHss9V
BF0rhWlGn2w4vSnvokSi8PkBCKlPN1rf+pnoQ/VvjHyz0JeJMkCKhPKwXbd0qJRUHbAol8J6C9sx
oLyQb0j4Y3WH+GVbPLtNrijp6MKERjvtS49utzu9f4gtmoH6BS4hnuyv7hKioRu080nHEbrEESso
bxeborXsOVBX8qXguVdf2xtDAn2UlWeCI/uOq6C1JYCjRLKtUf4cjmZ30Lvc3Lz7NNERTXC58vIr
0h9RtiJYsO4p6uj1dKJz8v0MsT4CjOTF+vuHjMRX+svd2Ue/eB7VotUB8Xa71+hPnFWLuXYV1UnE
EiVXAEUmgAx8B4o/BUBgUs35B/Fc5EcEHAo8hfXjyZ062ZDjPhS4s6O4HqKZVi5zFmEpIJJEe/Ki
Uu8K4rjzx1nrWhd6dXO1vBEs985xjeUM9S3RGLS9hnmxpc5uPnz0Cy+GGPZUJJpNuQH0qLBvKVHx
uAwRKxTU2WdAS/KR1IbO+zCOLes5ihPUpVUeIPa6h5qH4ga3H4xwAGmPtzHDUgoiL+YgxkWsOMJb
xFaUwkam41DF8dcCfOmeHcmrtDk7Ce7GxWmcC/UbayCXmy7geDsZCgTlmCOoo9xZr2S/UZxFzrA9
IV5hdN0id8cdeSnF+jWV7fwfWy0jOZmY+jmtqRGPdMRPhFuk0zRotjAdJolTLYJpgBADM7OuZEpv
7ZFG2m2TkPsQeEo82CDkdUnNQlbJ7MPuvDP2tJD7JTityHN8v98/Vf1KD9ZsROIdKVNwZdUqWDPC
wfUSk7erhQPgQDRO8JFCs1+vZhNMWgWPssPUOXtSNStO0K/c79CcqiEs2ZxGr1LsmiRAKtMJyABG
9ERDmwJUgF33G7dOjgNNjvgf0FXlMee2ykCYHe1bkwNAmh3aYC0/sJxGM5Nc2CXaDtoU7YGNUyxv
cStH7hJbmwW0HMea3yt6x0sanP04hVMxCIrjj6E5M7ynvc+0haiOxrxh1/6wjxfrhFXEdqIv+hmr
mwfZnD34xwLlxXH5Fodd1HgmJdLvbRdt0f/2bK82hA18BZ/GQ9y3AeHIqmBkwVEy9TuK1Xz29G9J
nTjsOWKH1ax/waNU+hv/WJmS2JzKHjj5fiekedHyRHTGht4cpvApZX7sHZcB5UEhTQE/sSBR8Lgy
U9OWb8HWCyKLstsxSol4vGTDCHOIBvvUoeqqXKa08nNaqY0lZOcKu05zG0rkSBbvs8U5VAuDhTnO
FOBaop3XGw2az5QKhEq3vKwQAucUpFp1jFVcG61YF1DX6dI7O+/kclpoJnRcG0JTHQXYMZvMtlIN
MMLJhX88K+AMMijpAWrlhGSZNRNAu+eRF13iypSaypXB+FdL3lxzF+U6uddgv9SpCEhtpSSxLL4Y
gfJEBn3PmZCSORSxFH/9e+jBg1Dx+XnFjwMBvSgGyjH0cKTLqpOZmfHg7QztAK52Hjj6tVS67W0O
v+9/Epk4+UiimgA7jw/SfanthGtmV0kUmZxhiwo4L0IJ7BsEPF1hsO2JZMXcZW+t6FZbPkHpUfhZ
dEEnQD3xRqAWpqmXUmOHAMSD8yS8U6sFqKBq3PLHb8pZtN6zFufeknjHntOiL+Xrk5ADgQ76NafL
3Vg/bAta8zKv1JMCARrHoXvIbgIVJe/UJ3ofReozi699vEfEfNKj1K8IYiMr+h/G/RvhmYl3UAiA
57XehSUSc3LgLjdy2wN8dbwGqmZDTXzBtSC47J3r6T/PQFEOi3Hxzy23XvvPQ1cZKpIpK0zKUBQ1
edRKxj/c+Zg7/9ZWb2WkvEruP5rR3ka2D9Fd6CRhi/Vl7RiLvB7YQgLuhlg/b20k9MNhU68TAEnf
nuGafiM8ikr6jvRbnCnWgCUcYD8oh1aRAYsIg+CdshUxiuDdlCEwDn28M0of4w69I4jZBuGv/8pi
p63J2BvQ9Xfkn5zA+n5MpZCeu4h9MekdSnfXCgnBsb1J4v2Nxg2biw7j3cCeErLeR5tMOSaH+D+9
X9pLZOXdiGxdDuy2dclhKf+V3H3Nj8iR836PN1nDwHJz8ucSpgF6l0LuLIDWz8vLk/3K0uWcG0p3
hgvK6WXWH7BtqFprwhq97x65kzHV2YrlhHlaLn9GgQjV2Zm5Cl3njMhcM8L5WyfERoHEw9AV53r8
p50Qave1DvSEagkl/zoenOKKKibznM7mMOKEcWaxGZWk0OMk3dRKnMiu3UnVJrHIbtSSGXLyZ8od
kg7C2moIRZa0jUcqtyJ/yUPZaurfUodtzQHYvSn1kMCEBMKlBE+o794mWYB0qOWUJMk9rxSt68Fx
onQtXNnewbioqtObL3NaUyXJQA64MS1LkIRE5U4ljfjClusfujlD1+x9EDmKqC0lrNAJ5/eaDVqV
wGvdRp5jdn/CfX+hFMBWzg0sT0sy0I675znuOPTOyFyQtXf50XwgOGQzPSAKjZusZtyAJVICllNp
pDSgPGd429UqQeTM0qepUarjH5egrSm5tFKyK6RH6PjLaJb0SBUfp3RLd9d1wlOaIEFlV5TMBv5Q
72JStXJgQy5s1dIKgIghsZd/qOW/PmBCpMkTlNzwLzFeZ+Gw5jmjCebWelKV91ctrZ+cNTsh6xU8
IlDOGzFWu+L/z+gGSmd/zqxV77iRtMoke450N3ABlDAvT+tlL2pRCF8zT9/Q1H/ePds4MILI1ts+
J6Sp6/Plhq1becrKOkUm8/ok1gzwblYzDh4LDq2iHDqObbZFu13QZrzgGAzKVjYhapyFzFEmSlis
yIVoveAJkT5LrcVnOkfu8sz/PQ64mZDvZBUrR2BTkbCJVwTK8o+KwlQ26z53H8Oit2ekjH0KXahc
4rfCI2528vG4fmq6Qg9ZjmTuFGONaAHP6YcC+tHk5P3i3psktB6u177IfEw0zz+n9YF7TByg/xLr
Mkq+aFD0vSngMp5CaugWqDkGNeGeOdqwIFS89UwLwZQ8y41E+1NJwgtm+ATOCetYJGjaGt2iOHl6
rhAjjT3wsOeBXFkhjOK1+C9pUZ9ai0zwWky5AgZZWnfvVit9q1Rw7LMJxIv9gJrz4dowdu8U5k80
ZAFmxSBqF2+xcHYRgKyzoCa4mpIt4GOBHEvBc7ne4D5Yzw+ZI8Ecf/VR/NEEbEXUPa32+TsxPwBu
p63CM697MCej/DBmGZWpYdeVjqCFRYy2dJJTmV9h7kLKZTUytrdDek25uHHpb9JPoRnbMKp2wf4M
4umZQpzzxWMlmseFhCnq0mbgMf5mQqmz00tcV0DBx7IQHL3oQkLj0oOrqsqOwZXlCqvJfStuDNKC
NX6d+WqXWxDnvPxVAkdQLZM3Y7Eyh3UJpUsZqxxT4yw/PzMUA2qD+DS2ig5ZecTi61z13vEcBlN5
Et9Gjq/6mUl5y1hCBvOiDi026LHG7QmoNJqnMhVgjeTGtR/ZMFc5RlHCrWifx0gF2nSkAD5SiJ+K
3toK88c48fqAsslZ1MHQl7Ey3a5C0wBZ1VDzlSpuClDUpdboKwQhVgiHaR4RiUKDLI1ed8l+NmqH
hD3hcDUhmdN15wa3ehKbJPA7z9WjxysfJN1pqvNt9L/xzCFkKw4xM7AMzpGz/of26VRg4BZy9mUT
OqJmUgjFOk8dsrc9trE+zcmelSm5l+5jKQxS8wPOTm0ju2MswaRVBLZq27uJ8hE6BK+9+8LODHxc
Eabnk4RpgrM3C69R2Y8W1wWBEGgs6J1I3v0ZnFddM/bQqyAX1DM0y5H7AvpjRtbqKfvpsRSORIx4
L/9broUQz/Yh9q52vR04ED81tBNjhRUDvovSQRbVlksKPDZU2gtkcJsyvNS8Y3RxjnE3VeF5Ca5d
06XnLaty4BKeEgIzjlDBuirFvG1uq5xsSqur7m4+y0WwfYeVJQ0eZEFUnzrLoeLHxg7htV9ysdcC
V4/1QWc4FdPNWc4SjCCmrEtmyge5bXFqaMR54I0z5okE3wvOVf0QRg48ppUwUzW2mBkLwMPuHniF
FfGZF0atTMSIZFZ5kkuRhl4ZP8oJj0kZ6DMnlS1ghWGrGX4FugZu69DfaY7dU/oB9yrh7QF7Bjce
UHNYHF11bmDFPurtNxH8gWoU+9qpYowgIetvQsp4ZsQX9+KEwKzz4RpVp6QvgxWR9qK3ywWK5np7
Xv/b3oYPAs0OjTr93wsJyE/cpZw87HV8C3+rm4MPGgQJeMJf5asfspcLnxrTdFyaqualJX4ELQjd
4BP2o3Tji51sWewiIVVnvF2RxCCyzOPU4MRlZU+DfrUFtRRMW6bUUXWsqGe/0zpO2e57YqoCb3cB
R4TAARDLZH73bFkHXtZaeZlnV8AFuvV4YLCnGo+Rf8PHvZMFj+vVPcjt/V6D4zp74pKRkjO8kAd1
J9bBIN5qdY7BNftnK8xzULvRbqChvpYkWMZaPPC4QRdVKsbpmc/JmrK9E3wR/6BVs0OdH5BCgMSd
ZnPnaI7Uo7JgbAmw2UameYCzZW9Du4T92yK/KMpRTFPJLrh1BI9lf08FaHnRTndsO91GZHm+whqV
MaAl7RQbm61Ko3rZ54qNB/xRzx6aYl3CFzllh4rUcnawKovVDYU5kxBGknmNrLb7u1hdCbT0TYgF
c80VpffjPF2PL3IalYk+R0jjzGJPl0HpKW0khTCB6Wlkvm0FfDF9HB3g4nGROlB9FwrBA0dtvc/h
XZRSg9MbuUuZ27ZPAvzDYVkgQjw2Tk7Kl1PnQLxOMHljkVXsVvd772LFOzg8AObeBkA0YY5fAn6A
00pkGo3ZygG0U4kLSmct/jajWqcrMBXuoWN7jGAvO3RkcjfRC7r1XgYVUXxTwhN+zfvd9e49b8PZ
vcRA7IwuGbZcfsRmQz5kmq95VhReY3BlJ6Sp8mLPfqAgshaTtDKKxsf6NayYO2iB89JDxBA8JLwv
Kie75B9FP6fryxOH2VImR+x9UxjxxOt5hmm6cht5qrVD9B2m+jzxjWuBEnHcU2MOcuxlf7hTYCSF
cGvr3R/lltyS9qTr9g+7JV1XQ/qjKuWVItK0F7BB9X9n783JtmOpsTZyvLEYvcjhlvGQ2wDnXjBH
y3l0R2SrfWJzoyWthXBAA39AAgd3I9qWuq2BXYGMTjrAMTadRbV6vCkz1JkL++SD/Zy5PyTHagdZ
aKQ//IPOEzXi909mpzK4SEDHM1fWuTsXhp81YJzVbIqXpPnJdU7mWUFeJmGCtYelKuvOtGBzqyAc
pfseIFdf6PQZj6lNNQPmH0FjhxA4+EyH285hSSQViswyRfdKAr306WmS03yzMXN2Rpd2+kPtEKNV
tOxVhFgkan/DMtuO0lJ3QXZkS3mzHLe+LB49pPa0Rhdb4Jmvng/rE/TuCPfsrKaKZzfMmfjqMGci
q3YIreC1so/O7cQny7J6GR8RmoUNz7Zqd8/hC1O8A0iJlWWA8KvBOSPc53c7Kvm6kUDFKDd9b2iC
jRJ/qmfhcaUtJYg6/JiOPIu6Mn/53gcqdj95MyZ489X3L/Ui2/f4nIx/2BHkRhOzWYZT2ZDefbRH
Hvba3tmyJXWKnuY1CQlY+3cF8QhFj/NPg/1pm+aExG9AIhTJVMlbylj8NzAaT/SZC5IA8O1w0Lgr
I5CHVJOPje+kJ6xLBe3NwkYmACRGpxk5kJ2/zhvLWgoFA3adTLb0CAntGNvSm4NcPOEmaA3JCjW2
teuFNL8SB9n5/C+/IgD1ycjqsFbb/0H9Vx+71EXVP2MjkaP9RVYe8ddsEB8KjgfUE/mpcBSDhe3c
4zZPFq2cNzYFby2AfyTFyGRd6hykzlLm0CcfdyO59sdEO5vLkZTfnbZU/niEucxcwOZ7O6yhIrmz
lXgS/lI/llT46Qt55xvQYRooP3gobrmaG6FgF1lYrC51T/ccbOIkZT9JXkG/bGJe5fyKFEaHSeQU
MTS5Yq3wpjqo1dS9aE1KXvrk6Nf31BVWBdvIUFsS6awXdLtHWH98X1o1UYlzz3rpzD/xE+pzlPoI
rR7pJ3K2i8ib4oZf7pN1U5Uuj51ban9ra8ia146QsqIUYveHsd6xTFE5G1DfyDxrKn3QcVYXP1h+
9BaSdqMeCtQG91ypyHEjj5/37/1Ytx/6R8itbtdzvQb7I/1KEKW5MhjqbwqLot7AUvVGQq8T7nIK
oayFJSZzUMEh6qJrY94y1snKqw8s+f1BBikPCDVpBWhEGXOFj/MJv6es9wdDiGLjZmltGBjx9FC+
ki+yZfvH1Ytes5cQsxgqv4oDfJsthw1nHbQ6rSiFFfATObFAMARqBgt832ESa0TVbSfG1XbXhCPV
871gje01hojaDhg9cbT54+DCF63ZYtW2FwqedraHyL/k5pO4CLhv1cxbKgoaMwN+XqET2CleWaVp
11/gslIOEwE79zVhISxrVpfx4UqZmecKcl3phtR95l0h9Gu17Vj2Lsk6hr/2kg3xtTMzoUk7HTnF
UTGUxNE/TCBPBfX8cwyEDxYaki+MWBRAjON44LqccXyI9crw70KxyhJ3cI7POpqf7kGLdg9Wuwc9
ud+bXPmvKnDuIoiM41u92uZFept4aep/80SHJWHG8l+bTM6CZ20Htk0IiW4JAXli0nl8EJKUIfHW
20zCbNdaQofCE+EbWl9+9o8NrkeaisSMHKbCXhQfbZSc9rCJABhN9MEvdgnU7CCwj+jqiWsSYhYm
y1W0d0HsWjqZVZcsJrwLzCnxjf3BGDup3K28lL2y70vSIoW3XKO3XMcQ6iGUa5dbd57S5kFVHs0J
iB5xhuMu1/zN+flbnk2iCpJaYN32d+WFj1P/JXxr03H6UmWfRV6O0qLve9T4cNbl/1+RElUxL4oZ
gkqF3eFJeFSupcXQsi8vkvv2gdjPzFkfYioPEdurSH6RyHqwhHVbI9eOll+kaZOapqBzsKqo3RCi
fdYsD5FzpFcueYXBZjUiPT5+1jczuD1HB7B74V4nY/OFp/zmqFz5++9KcIHpJhQdDe1vOFovxOH2
pmE1n5CVE98gvn+JnjbqjE5iAG/velUavQ8yP96v29DHQlrKIqfYG2MyP02HAASMQFgoeu05jSqh
wdRgij+IudF6Fj06pG41iezPiX6+BtQDiZFH/4qwEeEwwlsTyv2ntSYE9Hh3Xu/CrKriRqlxqmVQ
RzicWTgeeI36gUuqbQGbRg9FwSYscrgw0a5dX2TznsWR56h2Yrba6CLN+tABRfW5EsLlLbTXNpDK
ZRhYKZwX+svR2r3xrvWzJka8hH34BkkQgPTmSRBf1AiAebMgk4i5LMxCkMD2yVjl+N3QlQm86YbX
j2zoSPteKI6TuAbN10Yhim6g7tKMKJ17PTlLISx9NTn6RIAlYHNOYQoegNmKcBwtP26FDyfL/vSt
n20XPmrZFy002lEtaHgV6WKCX2qjnFF7I6ODtF6tqOWdupOVRS5lO3lBYTMvjpfkMeR5mm10w00g
x5lnVNb8iG56oJmBjmCz8qhmxWSsKRHahi19MM2bj00YEk3R5tYz4EYamFez3x0pa9nrQ55nEeFa
9+wuMsYu/iz1AMVXcm9lb4tTAkKwfjGaHD/D72gOqH/ziwP6cMW/AwYuZ8NjMjftJPqIqoquSGJT
mRhGqfk85Nj51GoXhX85khOJMhlcEmgH4CXXe2n0trOFI98I7GZBUecTZAs4URD+bhokQ+S+W5Ms
DSUXE4jGgfck38nHvmStrchwwDhM0yBxKI7KEPys/kyott9CVoSALHt5iR9AlELA1qiiiKLKd18D
cWV9EPnGfMxsX2WZqK7YnSoER8V4gKJcnt88W54o1S6bsdFk143TqZzpUR9VTbhGm7N/igghcHct
V2yUI5CaXTdENyKRwADMkuLYOQ5N8P+SqsYw19v+pqEQBFDl+0LK3HveVvU+gqAd1+xHNXbe5s9A
bTGKjLFelvKwUUAozIsP0FG9Axo7es70JKQTv+0cytsGDgN1xhpQLvgrEAYZTqgGlo3xVQw2q99u
3rG3WL1+bPjKwOYh2MllSJt/hLI7JqiV8SNbtzbJbJaCsyb51kcpofyvb/sIOp61R06XpilcTIfj
LKn+KLygnKJXUrGsqjTzbhzXMrWmgBwAWjE27pKFVFGoNQV+2i1NOeCpnSzqcS+UsntbATfsZWRb
nlTEKHOJM22HKx6+2QEQAYo55uvQg1/aqG5YYP/6blXshAkaLxswGPllkNZkLznvOX/2HSWTKS3U
X6tfroPBawYaAN1ijwSTmHFXv4Hvs2ayRobrDwpkGhEYggNih4stLdnAR5eqUxkCmdlBNlyMap6a
GhYZTiU49l5vFcew+QYXbyJ+aOO1yGMTi84mvH88vAPy/UVSJxn3GsUfPlBhly8eogXd/5NOQ8qB
6/lz01CesprC1ZhYlYEP7lBNo+Dz7/cdWttY0dfdaIXakwLlBvnq3xy1m3AfXPl+79OylJCWOYs9
Aj4v39tSsDRSFGpnqHvMnU7/0j/mKGiME9CJPfkqdODeIdw7GhGYagzR9vNhfM7cV8rSdHnjioAn
I5xBw0D6lZSIlbCwWKtwLJmsqjQgQcXRf69j9r8jMR4Pv/hlLaYW4c4V8MEuTOhbK8OcOk33wpOM
VJVi6F4dAlcraE8b+TgEqZPfZNXUrYrqSg6+J+RME3uC1ueNpXQqBrXa30w8BQD7tJLjJa/9Tpg0
1L/tPB66t7+Ky8sREMKSVp2izUjxvNMudB7m+B+3k/OMhmlmzzzPqF9PlW872cNRzuVMXIUyH7WE
zhlbkqzhpjKR4FdFjaG7mGO4hat4iYdSbzhpX7SvdiKqDDcAcg5cCX0/H4siRSD5cuptPyjgH2rl
piJW3yPKhiHy/rGtxZYV2oRkx/C96kPEMiNdVw6sN7n7KtzWS5OifNIzarRyNmUXWwN/85HYRr1M
p2uuNthmbu7sOcEhf3bEHlqUee+M4a0dSjdgYZKIu8Ra/6+GsSjp+ug6+2Bdq2VTwKuAlxEsh1my
wttGhSEqTwKZuT417jZmyQKagwmaha9zwBHZl6RSkGFOZTH9ps7v0oDKoI/joyDF4NiAzNu+EL/n
ALI1IUL76TvIIzzlOCS97r5I/h5dPADOlD7fGgYnxmrRSFbuTGYHq0J6QHJcNP4Fih9yUCDtQOIi
86w6DZ1wPWkA/4lvQj47fgxs5BrNVH9n9hABgnbjXIutqo3ZCgJsmt4l8V5apVhglhJG6itAOR5v
R6gVBUi6JQqkUF5pmNHLr+gmkYrW/UK70IZjkB6SvAJwqYQr+orcQ6liPEzuwZWmF+136bXxBYZq
na1hJIpdFU7j/9QkGXRwkHXQ9f7xDP3hVEgItdn/ZaFWcIkrV4W46ldieijPLLXOTgvbt20qwoPe
1raVJ4gIskJY1kv7ISEsTSvy78KI6zpI/ciE6pxo/HOBHR5AmDbaC4Tfr8TPtOV1+IgdJldP7PGm
fEK4RiQjWER0KLE+7aOoWciQy+93PiiV+NmdEOkntWZeW3w8hWAXMaExafXUGIwUdcWwRbhsFaap
t46TjhsM19MpNu6FOARGTTC/92NyzIz/6NG+u2YupyOW2Wa4iBuhTSCjy5q5X6cojrLvSQsihqSd
e6DV+SGQVmaUdI7JDXe3w4NilrmSOZhoHBGcyspyHQrwA6a67ngfwIbef3LhmqIKn9iOyvjQmyoJ
450yuT57e6BZ7YrmoY+BzxkmedWzN7YwzUG30eSK7MNt2uUQ3PCT+J2hIyt8EoYRVRNi3OtDbXE1
QxwdXg5mnexq+GmkiRoj4CmFa3HaW/QibKj8vKqEbdVVft/fk/sBb9tDV6AMtnBSldChETKRuslg
Mt4NX9GQabpIYhgpkHnbnCevnF49GjwbpQIjfRAgI416X/fdm4vKMWLneYex33AF8lSdRiHmQR3V
YWpkvbR7eIhdAW7EoleBbR0/XZmlbx1IQeQ6beKMV8U+eYQhB1lezhcoRpOaRSKWK1G1PW153V78
Co7o4f0Sabb4wwn1kBmgiOsIDzP8LkzEmGVHMaFpbxpBalKWJFU03TXzollKeFLsNec/kN86Fvzc
dPx6jT36DTYfkBOY4+4aW2Y/lkRmgEEMBmdM0ZD/TBDyRyDPiNJhEwqH4RN3LzWn3Spde3MOn87W
xr+j/uW8YUUwA5lCtTHw0SYFex8X2vICioeupdo3AVn03wzUhYyB+uRSBg1e5dQF/lg3+YhWWoHO
ViXyyHpP3uo22fZZH53wq5HU0xmQpy83TjdZQJTR04Ju9w+lRmZCoqb36A8SAn4y5QrGsS14VxQ0
rnhbGufdDe0CSSm6taW658svhQrFsRY4P8aMdFZ+B5cW7X4XKB21rq39h8kQg/Md6EhWBu7sh6TC
b8l9sn50P4MBS4Jhdp2bf+gyl7yqtHayMirABcoAn011y+bPXrwsE5hJOWvT8JAIH5PctYVXGakU
l1vGjmAKQfOr/j3MfISo+8Lw3oTKiIKFObCI02W09xzVWkOS0UywnxX7bTf7wWxtqPq0FC1O20bq
f+eVT7zFQ3PthCs7tDwXqGjn2oh/aZW4Pde9ZOqbZrVKirc7A+vU8w9jPSx6no3vj7gMJsr10lkC
84a+bxn2Vn8NelZAUZnc59UxeedDq1RqLFgx4BERmCWogXTf0nHjhtlcqOBZjl3yhw9cWz0tZuTk
L4Nq2lGOvomSgausird4RyaDEjYE7V31UcYDi7SwekpN8dB7XPGVhj7/vMTl29Og+bTrTwfGH5g3
p/R7n85sdYhhr2EUgNniu3+mmcMaCUgYKRpbcx1R1MKrrakrEoIRT+s/684PRaadHJJWZEauvNai
91tCuM5f+iRufYJRERc3aV1M/0vND01izsn9YsDWeIKCPDtzhZDrWO5TvXwyFAagg2zpFGK4J9JE
VLPfo0qcWKkI6aDlNVN6cHJ6X3E+DLkcugHizGIZlqHkQETaKLK7BWyLn5xC9+GA+RgnEY34SyLi
1wLDszRmjj8UDd9zQFbEAEeaotZBENl0STGz4xveJfgyUqUaME7TE3Dugd81q/XDJoL8FChuOV8f
RWjIk4vztQt13FkFxDSfK0RISdTwrSKm4BYg9KPc8YMkkd56XDTsp83Ri47l3/06dhBh94NOGAx9
Gn8sWnd42fOIjcSnSHT262KaOyb449/johVuY43KFNLGndAqcx6OUHbrV75I7WWiXBhVy5Ma6jO1
0ONPoFoJSQ7qkwD8yHhF4mNsBDIWChx9EYwTgOuqfpKyJ7gIe1hDSO12YOI8EPy9Nu8qdtp8b9Hu
k6UJgpBQ48btFJ4wJ+kF+bd5pIlFLreMJ2EtYj3s7sKore/McXL0mru35dWRuZ0XinnnDLvzFbs0
Sjv8wkURaAGI9uWucSNu3GL39KJQgb05F/Pkc1DQjhpfRXBTv3uYSV39L1WAPDs2zUDzJBhlU7mf
6smViadhV6KscU5aB1/+lb4SHBQGBbqQTMOXBo2JShle9F0tCPKTZHv3dOYO7o8DxHorhNosUS/7
qMOsbQHEsm2KPxIH7H7befMJmr9S8hB2H0q0BRY0yTyz4QqxyTqhIfA8HuUB7DZ3/S9eJD8AXhmM
6Pax8tIL97eheBBx1ADwnoscoC2fqXv6EcsWF/LFI2f24UW8SrKD4Ra3asRaSLqr/taXaOLcGp3Q
Em9IiJ+J3TDf9ElDhWLz2MDLcsM877UtwLpu3sYrmMMPtdnO7+Q1MkXh5/aNL5HBKyI/CfSsUEjL
lLHrZX4l1af1YUC8YieVXhj6Erf3XA6RY5tqutoSEnyWOLZ8p+vYyOcsUQtx9jLO18nkO8oBt4po
F/GmJ/u6hYZ0qjytqK3EVXWqQwMGjXyClDsNuaRuCb4FgLFuOhTImE4BqzeTt+wGJae9crSnTPMu
s3bgrh596hIDlPftYVKeR32cCK3aJ2ZjH2VsVTyRo998S9IqNv5qOyuhBPCOuOUojqI9jnOaB06i
CTWQkn8WCSUuesKVukMmpus7AkzRvxgCvWi8o1wOSDBWoHPI9eU29d2/Bgy+TKhG0rmsXW723/fk
L+aoAgnov5Okt7DXJEMNdSyJzo4G/Shh7BGyL1RvLMNlz+JCukJ8JgE8S1+CucoSWiYLr094H01L
YHE0LXZQmlBogLQnJtIoAh2w+FFrexe2tMCrGhaOVVhY9VFxfWXWvpuaHqBuUxRpJBEVUy1r5S5x
gfRXMDO183bWXZLWEUu7Atolw5kaBQtR3ZxDI7vtBxtZ6O0Ph/UcspI3uFWZqAiyQXzpEBQdwuKf
knFDExHz5DLRAReiM3PetWhWPIBkIDjwoQJDOg5S0XSuTnZraG1znnlsKhukNsK0Z95pED0hnLcF
aF6dhikiBsAvPYktS9xMHIbth6NnySk1QJYBTQfzuHMN0jAT6uflv4Y0XS/ngHYp2Of8AbyeF8pJ
R+J2shMmh9mST277U3TXdKby9gT0nwucarSZSWbymPGIc4+A7A6KdQgH/TPW8ZbogyCqzpfaKGSJ
0K7/vqFAhmG2LLtIYVSwVVe7rAuR1sZkPcy8hDBZ5BPFJcbDmcBErLyCxYE84o2vzXzFo7nw1Yo/
egHcLJLuANOkK0FwCuNA0xnvxU/UGFgnpGpQxXx7CrwPgLPLycYx5f+EZx+bStEHYBhvNulFEMbw
w2egoSDRJDhAXf5M154gA67Q/p3IrkHCBhjSNWA12Ewbatotovt9Yp+MuYx6EDxYgCRbTD3XJT98
GNnvufNRBuyvGMNzTf9J0dzUk478YbHI/lHz6Gjle/CFr026qtH8iTHjxMJy1ywv5lhxDtarw7+0
tUk2dhlakiwnsBU6iZr89BXIU2C2+lj6lqJNt8AsG7W0PhVe5f5GOZK8lCW5X9Mw7nKAqEXBZgy+
ZbVIDzcIXc99Kokcx6h9qvW6oCHDBh9ji5hmQwqlTPx5oQv+NTyBp3Uf+Ht3z2V/OunUey9nmrzs
I6x9BFBLTAbHs35YVlItsxsJAjX3Gc/EOl58qGKHdsRkX81xDCe7nt+TJZlpBAzOk+YkhDgNX24r
TvXwT0JK0R4NZkzZ/Io3QSD1YaSLJcAE9EnCgftD4VQBG8sZDlMbLmW1LzDix5H9jCFTlnjJLK4I
sqUJt6/qunVgwP624i1xEdgh7K8uRXMwGOCInPQtv4lVVlyr3iO3c9PZRYSAhQh3uG6W4UcCUT7C
CStVEhpsG2D84J7Munj503Zs65zc6sPgsNwbG07zXv8kT3l/3u7Tt5zu9IW4OlEtsRUEm9Nwq9dc
slaeQqdj8JrwW3K915efdYfoYDto2vCTA+HVdcZ8n+BufuN3CS5Ud75VDsi+ovJPR+6Lri3hVpdf
7ToediygIH6tofRzYCwivmVTaImUE3nfkrY053/WPzucAv3tUGzWBjxYHN8Na8xJ6FjVinVnqEv/
h4pdtVG96n+ZfXCzlkrGe0g9IgSMpHmKruTd46CAlZAQ8iS3mRri9OrnOh39tz278f0w1WvRyzv7
3OD8VoKSbFYO+lVhZ9Xg10Gu4QBOobgRZdftweCvGQNL/Z6/jz62fnzI5Lfm0Y7wBLPho5mX0G6E
GgUY3PZ7QYxThdjIvrd4ESfUbwM98PeI3N8SVqNneb4TVv6YRX/4qM4SuEXtYlKW+i1e6+tvuHg0
2nh5uFQL/q1adM82LD/MvUE8RnTAajbeJcB1LzuMt+rUzLHLGWRTK1WZBOmoPSTK5Oe+sQ0yT3og
MRKlruSSECHF39bfHb+2ualikcCViUHsdAQ3RCFp4QycyWNgMjaSZmEA97iYG78YsFQxFdNxPQld
OxgiA3BMjlaeWUun4Dmu8P8xvXcSQpI8zPs9JoiyD1edKKEc2FhYy/m1RfmiM4olDmLTS4p4auW1
AC7Ub36OoRvQEBVe2h5fXhfDzFHS5CglD+NQivzHHoVSCaWjTXiU55oeXGtBFD7BPLYidrKvH4+j
Asi82mejlsOwaXSYBPobgQSoYLsVmE3g3yUMTM/wwyyX0xKhTz1xhZ4uwAalu3rsovTKVG+mXXhq
bzZkMALoj+QJi9hvm6k/Wec3tiI4DeJfb/+ipjsuXTsdIGkgHGP9/aI0nqUZijeDnRzEZi8SmGzm
0TLw0ELvEKmAYXP1+AHl4NLDjviNFN68um3eysghv03kcrp8vEh7jnRgXSjv4Rkh4ga9AoJcR/KA
j1cilW4YkUknB6xxqp/Ny4Lb8C0WMJ565ogMPPbX8UctRizut1CGqSfrzmpHLd3sfj31YcsR+aF9
HuzCHUh9jWp3mSIJRrAh4e3Knkk8Eab4K9O7MbeIDI0Ls0ujx2SuupBgOLxJbOkKhY9pdDP5+4DT
cIOjLOErNguplxOxpkImA0EwKSpzCBntVaf+5FTE3omdqqUmws7l0ThyXvbYczTrCBhd3ab/yLCL
mlgZsG2hJeAk3JDHt1bo1Z5FWln9DBIiPMT948SNH/USk2NahvKnJoj6OHwcmtXZKlaCchS6cdTU
t7g13mkG442N1e3DKOuhvsUamQiXW5B9uIpUrupCK2uEDblv/7PatOjLfCaf+qVLrix+ud4oIMvG
p8O4rjUUkHoUEf3Eqve0cYOmr6A/TaM0HTv9yCPCDRMJD/nnKGmsxW1Eyt5B0KbmNF5A/NazF3iz
njWvS0owhv9axvb0sdUaIDx0I7J8u8BEZ7SIdvJ/GVZG754dtN1BA4iO1MVeSZ5oiJTLIWUP85ce
wum/zFXgUKkkHcOZVFn+MG3QQ+/PrLOEze7eM56+aRX7RSArHFgaW/ickgLm5+5//5OiwCRL2a9D
6EKls5RCdVtoSi/7S0RTNUSnl4rYV6cYTIzYRoL8VDV29uhrYKWs7v16lO1rkFsQz5baLH9Ujx2W
HRe6pBRHvnJbNVs9xXRHWCI0qtDH0KOVCvQqxuyvV3Mq7RIGw7shphCnjYvi4SFACxqwX1q4/Llb
NqM7AGCaciJbnUeZKCPyR5C48R3GKLGr/BjzQVp0whGcvDZ2NPAmJpycMDqJChkQi4j0jHzDajsI
WTN+xfKUZ/rzwzSliHgf2pn+Z2LHww4cwRhun673YzkOJAOA2G1TlpFTSbTpS+vgCAJlrt7RlEnS
ZZzhe83MqHOSvIPBc0BobxJr68vB5XZNjUtQEC7ITs9eSF8LrlQdhhsxP14tsGR8S4SuFo37A/P1
xwtQfvrM+vzQhI/Sr7oohh80NJSpHx7p/a6HL2F94xLj1byexvP0lFVThIujmzey2dIFA3O0LKNO
xlCTONmWJNyQi1T5HPd/KqV1xnplXRGnxfYsjlPi9QBKnNf6P9bnhNf5iHm8zM32A/esGBhNh1oK
4Z0xz0fGIqb+p9LocOi0iU/tAPnm94ETLDeSCi8aocavsq/lBFIlIpJscpYjQO2k5PV1jzOdYTR2
HbGMdRRfQ2Jz5D5HRedm1H10TGdwJ8SlvUI/PyQKUy3F4dSuAVjUAK8QTAKXOfmRqoUaqLW8XyqC
SuwinflrMVHtDuJyOj70B/L1K8lxZ7AaQP3O5wK8pGBwt0dU+qF5J9dxrzqignciI6LmVxOhocrK
p5rDJCoXyMwDFH3sOVVHZXC3/q7Nyu4PuH2JnEQ4tSxR50nm6yjhxygsEWQz0U+Vk1k9yeklMkRi
4duY3YL/3qJ1fq1YVOE33x+rqOdRdcLByg2IsAgB3j0kDN5goum6jVvnFBMlrHaBxcfsEAmQAHxe
H5HSDMM3+xbfAt8fq6GbsBvzytIhEcWzaETM4my1769Sj3//22TRDrNseuvBbTova9YTO8XsQ0M2
yI1nv+wcrtk9MnTygT2REQ5Ez2osYy6dX1CPA+SGAFKwsKrIn0rozgkK9UBJ2/skkuYt0712Qpco
Dware66wxJl8+J+90P4Jgq3IwyBXAVxU/myxU4ObDvcRP6UXgV5hzARGn4FQDs3lboYJPB2Bbt+A
en2yfS6BVrMqaVlF7S+qH3zAkunvkQVOtlizTg1G5Fu+nM43f8eDfWTiw2rWi4S+TBabpg6ET+34
vzR9ohjWHwv+2/tPX5YRnVFx5dqyS9zz8Mi8cU+7qs8bl8VIS1gN6lJTDi99uyJFm4c7f8DSv7cr
1BgiY5rP4oHtx6Ss1myQWeZ8kQgtPxdbFU/ysYX+Dhc4czXJ8ux0KILuF0xj/1Bb8v9P9iL513kZ
G3OaWTcriK/Jh6jmM+8eUFZrxoRGNo7vsSfAx8k/8AIN9exc4S3UhcJGyQXOn4zof3fVTunVeC1U
HBBeo7c+wG0Y7EzvxY0zrxcCDzztfgpZGJRMIs8Uy0BNqS1hoVJj+U2N+celHVNDzEJiethEuYjc
LiIb81ImxCoNVFjwIHykhwEeLLCIckfOWyX2Hv+cFRV7fkyxgFLzGPNP6XngOrBBlzl8bGk851hx
fCbkawyJg52HS0scPmBlxJCCfNi7lHWtC7gKdoUHHh7VGHi++0LDZdSXgt9DP7S6FLoS++O/6KXc
9V5uxV4a2MBYYqdSDGT+t616TEMZLovLZuZQr7dxgYl+bXeqLYWIPKwRSthGLGRfn/HDGaa5i5o5
QwK+8fzckoWj9OFaTkPSneafKKhH+rRu1hCgC2G5LjDXVNPjCCnMVQNsmav7+fdmVnV7HS+A3jkl
G6hfwwv7Mo/9U3TPYcrHHOvVJfJKn5Y6V2LA7d1oJHcJ1qANpidgaw8tfS4b0VMwIACKSJK/dpux
HzE82CW3p0f8h5fcnPXcAJk1RWvv6Y56yLMMdTXr73zuOKrPso51o2D5oHBuOrgFhDm8kpgC3lIQ
ZY7zQ+jQB+3Z66kvMm6O3AZMdRsr7gmFMeixtM7uWAETUWpBIhIW/coJVTnh9JsaGnx/2gsngyk6
kvFlT39qYsACgGxFru7WFH3NKCEw/kxGD87jCNY4x+pJnLJjz8KZzQw2jCfeayMvLk/SaKRo3yd8
qmK+1rw/GzJjRgW2th9hf6pTQeni3tjwwk5MntGP8eULApqI1EzMQzTShvxrPnyCEuaAGa2Eokuc
ccWnabYH7bPGm9x9zWDJcvlhdlfTcuj+6uZPpVifCU64gjU2QEBdxMckztRI7mDyqcccREBjX+7N
siRT4lDwaKl4KO8pw06sQTAOpLtCJAaxT1UVvbEJZzzqqZsSbaCLSIfL4NKu0fauwP1hhNaBj9Ji
53xxpt301jqSZAYddN+VDsNGw2Epf8JOpLk5Zo9VYYmD9oyIrIeH9JI1TylToDn0zo8m2KaCnhVv
hM04yP12LgO2jO9WGOxK6r7ZQZt1m/ih4dBCDQbz54BI0IPgJ+D8A8/hAGCI0CZUD/TXmiYrrPp6
ytT4KUr4jdo90Vd4AaeGa1jV0NdZ8AaT3j3NBgJzPpNeJ32Q8EzJ7Je6aXvsD8fuAZF1HSG77n5w
pUhC7AfWXirAL8JPIvGEHgsFXegSkQzll7Z+oSt8n8tAC8NoWLL8vns0UXcFjXi+9lRr74Bh05pR
OZD60YL74l+e5SvAiXNEItUswO3W+siWG4cQ25kCqeDMorXaNQcXnw7ddrMqVj3jiMotSIL7yYV7
VyfhwYC8r2MF5CvGx+Xm23bSfJdlxOXNpVSf52aaCRlwarPGWhwEc7DQgyrk3U9/LHgZ4JUg9+Vb
+BNbVFARot0Aodkrh1vylw0PoHMDGZsnn+C5IlPmYZ9eOPhK2XXd+/qFXb/wiVSddLH+fbHBTeAT
mQolXrtA7RX02XNMiWOL/cgHMS1sCjTG9L5DOtox23zJ8UdSvjNEmLP1vZSm1FFXuFOp74rcTkgQ
KR6E9L1+k+X0szFpqdT+7ETIYMYR8GwYY5rC0Od0ehS2KpIAGtt4lGsJLe0bc1dh6pMM0iDWbVL7
NHUh8/JH4z+g93fWK/SHPc+3vuBl7DWisMi3TCZQ2/koo6QfNlUsy1tAh79ZLhSb8/L7cj+eSaEw
RAMFyfape3aWnr5BKVv7udCbZ01lUqWBmc2gGxOrvSyxiAQGBK28OK3fFRC4UxfROGd5rUU0G04Z
YNI/NMADycTJX3IBO78A//Z7nFtsq5BO7Y/aq+lCc7HrtT/ZNdVdcohJpMV6hH8QKzlipxPrcszX
8jw1BsHorj79VYjVTUBUvMBNfXK0gZUWo05WdkhdoNjGWfFq4TEeO93ygGKW7TxqJMRFNkn2BeaC
UZvzKdovY3eVNzVnvHAWJ4AqA6ZqX9jI3CYGzDrso7fJs/5kaFaOtOJTRkYV+F5NhCdG3xI/ffaV
O8Gep+4aWhS6YMfAqG2TkKnWYnJ8b3QtQsZnQAePlhNtqe1JQafLncTEFPFMRaZp8Mbb0gdJDAdb
NSUBBpHgMw+rjTD2k21LM9YXFLtpgXWMceKIklYN3BLhiZQSlGKrBjTYPZ8X3Nemffy/efGAndba
GJb1l3vEmwEDaPE/7Sag7AMXnE5VprcCKtQPxuzlZ781Oi1hpRbfphBWzoWMtZ1FcWSI52Rx2qnU
XjVnQSDJ5Ti6kwU6/WS2x7MG6fYLmUZAS0ZaPBGLr0thjcWdvwQM4mM5aiQwmaEulzyVR6IOzBjy
/QtRrU9unp6lQ2xv04VDDymoQex6SH5joTtpVZNFv2eeN643PJrOaNdOanshP3TGH6pHia0slX0z
StIEgBbD24b2DLV8hFm3tUDdRosEQBJeSf1EAnqwLN6fhKOiPP3cUvI1MKYhPqO5fw8PMSUYNJmY
QCgCA+0YP1NwE4XO3iBcckZXUtZfuHh65AqN45D2VGWU9OfPv6vKnJv5PdBxyJbiBAcohALV3nnG
MyTvfEhkrStmbZEnbVzHHt5b9t95AMvb+4T3Q7ffj2VZnQY9CRJyBzthuz3KvKlC3O8F1rdR+b31
/4rncx7Wzpk0DqCvPWnWABVSldmOHUS7kDGs+UyPBe5Ho+H3QX/Lr2L+l1kR6krHQ3MIOsczgMNe
BH/w4LvXUrggoXjjhj7Lqu0vb7P7CGaV96hQ4ScTJS5oT7EW0HgyhDukD3JaEZiOg7cfBnpW1B4q
W6TbqmCF3ic8td7AVv+xL514oQPJqpQnuYdghCUC6U6a/ZkQaPjbciFFBS1ceQKXfgR29H+4rjJy
Ooa2EeI52A+DXqXLWKkEFoZNOpCLrZhrF06JTH7AlDvi74mxuqmp7cu08/6+k3GNmz853j4sABzb
GYEcab0Y/y8/YPHuhVobsvde5j62QxHQihQ2jc1ziKkti7vYBb75s/44FZpJSrcgz72Ra/dyHrxV
jmmHq20lsZ5rHw0zCmLsCIwMiC1kRxa6RBAg8V03S14NkJTHsGQRWH9QYumtjQ9gxN25Wc0sYUrx
0XQkrz6CEFpLrcY1EWhFT9K3D6710b0WqjzG4ExC+TUX3hmNiGP+vtckWojC9s112xt8JAgKg2n/
QO0w0BIoyNaDTFpkTOIqvOOnDTjZn/Hm/2u6kLRVNEuV6l7fpJ8jz3CC5+alQrZzELzgqmyEOfjK
7fskz1Pwa3RQHHsYMAhb8rH0n0+ntmFfMW+9PwOFwQjsNa1R2sm7kyFfUUSi7VJBKLbSZXyYcF8f
gupV39UeGpwbQbMQv2+cI6idBShoKDVsTqZk1CNLE37Q6tEtaC5elgziw9hbKgrOFv+fMdB7T8Hu
ldU+WQyQ7uG2ehjsRsHKPRSBUfyTQmoFYy6cYLh8LQ66qK6wxNNou3OEElFTzfQNmcvtHawUOtXp
AJMmqb5yv7xveDG1h+3BUn1luyngTIBnWu6dsmpO504mSK2bPJychyN59IA2TiCXrMm+MV9nKk3p
nMtN+c1lHoh1feQGlJvC4pzp9UI55Hzxzveyfs+s/aA2cLA3P9tOKjEcNCy0qmuFO9bBqD88koaR
g1RQ+eeaSnHXsbbNXMgTQYVxm2fY8CIv0wYRvA9TvQ0KC8Mlz+izmx+IQFRwvK+XrHUkRtnI1kCz
EO7riheDHRAeDRJ6TGHwieIFwLGgE+WnuUFeDuT6sXj45RVV8j6afucKf+SVbm3I6p0ANJOBqHYc
mpRrU9Ai6xeiG6pV80tveMl+BlVOrsG5h4j5qlSuN+XdwCdSLfxQ7j6Bxz7FBYIhySutnEb8ZODu
DD0MKBPL1BIez14Ow+44yMp5KEATYxZd0iEdZIRxFNzkuUk2tTp2Jydt+HxABZVR0YSnwtNZ446c
CxrBvNkT4UzT7z47cFWLlyL/pwKk4CVVVcBXGfQNLypsBHW4rojuXGP/5bNyYSrTrjaLcay+FY0Z
l1dHusauLOsHaPqKeReI74BDnz82KcpQXBu2b6QovCux8E2iRlk/X9ZJjYcU3MCpxlMQ4xvgCUTa
gZJ6xrlvNfuLsmx8P4A7TMFnqWwzL5v8YIfq5+TvgANu31Xkgg7SvvS1i+chdFef1fHvS1oVwjN7
Vf8zFvNvF+tAzuvGKHR42MSefhd8eYZcvxuN3+i046HZHTC2QyyfNHx39VqWIpLWYe9la216CFYL
LiH+GzUqxS/Ai3xiUMzBgjlIVHXBXCfZIp9gIdIf3dSadL8PtWICVeTA8f9gxZeMuX9ILFKyTVLO
lRjWzDK/RB8cPgUGOkIetZkEJxlxjPy/AfbYNTlVERFjsJMTI8MFOmOlmA+tt3JmDDsSqqlJHUun
xyeaTTfUf6bO3XMbJhb+DX406YM2oekq4mFIr5Acjf1ga1CjHc8kzOHsk+GjmVWo4HKJfHDgtJA1
ngKFpl0JeLpL/tq1EK7YAidgO/DsWSj2CrOvAkwdjbsIDbXZGvRYbM4m9EYWBfX8LE1stnYh0Rg4
zJ5x46hLtdoid7KvH7iMWsYnIAGRqiJwWRO5OUAntZXCMrQ9mu66sOtueCTVDEkNVCUFVoq1xrSK
91A+V2CXUwEXOa/D6UF/u1kXnscHh2NgCJcypXmyHxtkohfmeiktFB02iU9mA6dyThP2z8BK6O37
tjj1a8Z1a38MJly4tW16qT71GUuLRyfjMzjwYfKSiFJ0hSfa6BKnEUBsyQWVzrqtFNfrspSboYRL
D0nlGMZ39W+iasaZa3ttK4XFD/LXQ5tNS+/0wNilLgw+Ys9+k7GSZt3wId5yeU+kZWFLuhKlYxhv
0YtbcdpS2ItDQpPIg/IrNkm0PXFKqKUUGVvf90vk2OP267nr+n9mU8LTls0zb9AzjnV7ryTE21gN
rP6L5xMKWuogxpT3DZiWeaoMCr3Bf9kRRTmiYvZeJ/RwFhODIeeZ7MaAJHa9EoOND6AC8yRHujk4
sCyoTIdsfLX7W+zwAfFljS8IYhl4QdMbmVV/rU8q/rEls8Zp2c3SXIUmgEKm3vwwjmbbVghoIK1K
FNTBTQUarT19Vn54fdZpLyLaxihQMsYLs27dpdJq3F7qEzZFiBzMGDgdAbyFCMODR3udguVSZ2aa
cSct93+JEQQrz+gQHsqPGCeNgQ5/ZVhgb0A9ZQ6aPLoDUP1KlcU2l/71sexr67oxOIO3JjDLF9cB
cgDO9ORzp8cXJeBpylrV3M2dGFfkqMjJnP8sk0OQr/qzQuF/0btv/jzszXdIbmpqvU0z2Cel5lrr
O9Afx4TDIg+ym4lPMS7OXnNffa18Wh9TmrgEYAD1nDo1tnkDz0L6/XwIayQ2+C8y26rJsoVu757C
gkyAnoIv8Si+ba3gHTksSErxLNp+rILDcz2bVEy0wNJRej+0EYq6hXnBe3NUp5wDOU8MVmPL7E3Y
VOx5vaReQL3maRh/PoY25Sq8LJZwjNte0Ivz21SYesWC3MqU4oPM8y/pi+6vzIS3NZ2927lIt0HP
UWq2pdzr2PyX+TO+FGvDlLKGFljX12hCOrjvNYvTIX+bjtrMy65Pw6pGeHm+HBsCIGl724nluSoq
CH6WOnW8Z1HKb7o/2uR59JR2XX1wjKIP9TBC/+W+iy6sNSmfbXmt6jkaDWFoLl/kqDczFJeN9HRg
zmsiY9P1rL1YsgH7owf6qa+vPG7rtXplGxSIx6x6Jf2vKV82a01uCfEbNOClwc1HyO4AKdyyAjsw
p1KDrAoe/IN+ycPPVo3T9N2K2Qu59ZrEEKIQWBHkccjhbAZD3i1JJA5JAbZIb270XkQpVKDJZuJu
Ia2jGO5SmM3GqbRMyvdYbKe20jEYB4mWH25mPiorokynxECTlEDbsFvtSMwQk+afzaiv+zmuFmfS
uUubvYW5QarTIZPElBaqdNjr2gvK4xLvNcWJcRxpfRvNTl59K2upXIf8azLvgJcLEV/1Bsfe88Ip
V4a6I1dRsT+7zG1/lOn55ShorZ/n8uXG2eV57BjmcErDhU5j6/7ymkH6ovo3qciH0gw3tCip+i9p
gpnJgh0UtovOyr4TE2DDH07tTM81YS7ctK+qB/njUeGxtD8fcehpLB2nLaCQNa9LZM+SpE+ZlvZk
RuaiYhaFP25i2ZIeuJ06puBrV6CHyecu5To1zncuailJuLI3fTnsstqmnrjj9YFMjO3DVRwbBG3Q
cznGiqDc+KRnvtebyZnQ85BQDWALZO0AG9Sc6sjxoqbatV9S0BdTuLdHYljyWDMRwRwWcJziTdvt
WaONhiGcHL71YJCzf3Ahri9XwEvb+PxOxgzXwAQy2Xn9xgsE2DUQ06dcxiUuQhUt89Jd8ocBuRDz
IESFCWNGixldCGvMu2D8rM0RHUjR90QSC19BtWyKWXHvf3P1eow+CrX9jbto7gZnzBfOmsgXD1QH
F7MdgozlNeSBtUFTbhnql49qGnzJfXKCN1fl7cBAEiBNPh4t495qmv6GXXP8L3Qo47qTLAfXaKnY
C+Qd8UMMoOPXjFJfPGlrR/stk10+eawbx6USVxSMyli6rw2RLvAwiCE2Z6XLiDR1Tb1WKFhsqtky
sjfjMTbEFOwx/TgHzV0DJG4Dhdeh1fyh+EQLgPsef9y0wEuwA9QErHFPdjeKQ9lVWmaE8CNCFE4D
aeOhboCuYO37cVMBjIlPN5L9RxgWjZt0uSKYiRufHc0P5NPZDHlLFND01BmG1EdGboXTiaV2u9H5
HgL1RToZhPJl8qXvcLzkvF4SrBBUx0Xn2syoCd8YPXQ4xZW7vIsFj66wY4ne8OUIJ8gNGeEb2Jx0
/nw2KxNfXmb7MiE/jA/p6TeWcB9OxbsE1yTjvZtI030YwHqsng/uVpIxDxSuANOX5Jy+vJabv+2d
LUsggLm1W9P9wbmdTLp1Sv5Ed7jH+GUSyteP0sbNq4MtB8/wiOSXeTPNMi3GkEClYT6z/qcXzY9L
3/dEBfglqTP3a6L5B5kdb3MspxPGrFWZhkrraJ6sziNTcp+vy4pssDIiEkIVODtDsx1nJKHCkrOA
gTBi7SmiWE/G773EAND386IaveA0zB+oufsp6xSXApPu4NhtlhjuZpWtg0irXhIgTNRQHrCGvg5+
eyn7C/hCdCVYSuyaTzM0o9lulG+prXNBXndLSkbLu5Q2yc6luFw0/gbGNYgCD1iwn1kuX/933oNQ
sj0GNSyywzlP8KJpeKshT9Th7A1OdboUer+EAyY5ZJ5qHDdXiVVlg1wzt8cg98nyS16aoW8/Hhnj
jOk47MTnTn9mvHIJF181BWzjs2nIRh///qHPRM2kabmIP03MCFNtJxfmE1ny/BjX96Jsv2CgpDLI
D7AcnoUcG7W868GVJgWYp8FoG0+xqU6UrzdbWcw0iqJoi4HfSWfoQnEKj/EvTtMI/sFXbgXfMqfh
g2zeFP0ePjq4aman0IAEtmeeOv8YdCXVZEXo+m+i0ru/DidgQYZvDoeRv73KtERJsuELvId6+vD6
BqzzjpJd3gEtHSI3HvDADjNsW+sSglpN8xLyyAYjoYtHaksr5bkKP4qva7voqTDbYNAC4mQcSz3f
zt7GT7lzc8sEKQ39XXQqwtEocwO5hDtWfWeoaloT1bF+GN4KrCkrFawThiB+UKT2CYbAXU9aRHcn
oCpj6xjBklqAP54+2SPzuUytT8V4Mn7ltK4omPhX82bJ0fYeJ/mxb2SJgZSDNTIQY/M9Kfl2/PGA
Hd3Obbbne41RQ41rkV5v77vW8vpU6qdtHp+djh5OWRBR8wCRJZE8nufBFEcImzZ+qwWEK5SqGecc
T8cIu6NUDUIYqzFta884yO7m4eMLPfs0JuY/SzluFJiN92kkqTzz7WeAI4H56bp81lNsznZfoM11
l4XxJVwte7/EoKmhFQAIbUulkfzbMLvCkssVlH61y4KmqvWHD3gtPF0FpLQJONO0uneqk1HguANV
d9lig9881y5W2PQ3caAWwUG1rLLiKU4TFGh+1pVfo/7cmrJqKcZlVXlNmywTylFNuD0mnGDmX6iq
Nt32vIvK71r2feIeHpDMzLZvpuxJghDA+FhRNnH3bzfb7UtkWL//A6kFYuouawC73W2Zlh/y1eNS
El+TNNKwz8lVex7o5oOo4217UjGcN+Z+UlEQibLU0mUxPOZxVQk9gsXp1NkR9OMVEb4TYmu/s6GO
k7/y8CZRpF480S6dF6bAxlmrNrCInjcxfY10v/q0aDMt0AP+xWZGSf5X5f6tOOQckvPTwP0peWRN
ilR40c9ozIYN6spOdHuoTjDvAV0iYVhmGKJetHUoMKWTmNGYhkXmGp6Fh7RwwBHnPPthi3bX1xJ8
gmbBUwjo/V4oRD/IvwPZDpiHn8dDWviVVMkaCkbsHbIWGDnG7BA1OgPsNKkZ1ZC2pW6FaeSmyYWH
RA3rguatYx7DEOTdRmFSu3Fr2A7/N43/MBVoNQXeSFX475WPaC/LYnm01uKhAZ1KIb5MuvIZWPN+
HRXW4ckPikroZc8x6X3NwNI1AhhrQmHhyKRx9sCSakZg19c3uD1ClaOwXGaWMO1zfKqXrIR+G2VQ
hiBmv4v3ZgwJyzbBUtDdgCI9gWEmcVPMo4bJuLtXnnyBFDY30aAjWnUe4X0OcZXMr9mYbaYZ5xEr
EQulgnPvFBgb4c195OHIweznTK7eBGu9ST6+eTMC+h9xtpTXWPgdpg2/tZQFRJKzb4tNTQ1yT6gR
3JA6H956ScPcOUIkCSDOroszQQEbnSevI6QQ6P9CTAFdRJvw/CFJbMuJzj2daAVtCQaC3HQBA0j/
iC11H+l4A0ilXBdl1/cL/OxyBsB+H8eOZ7eSDGli213xNIErowKUiEInzUnv3hH/hLyx89qCaj+1
7Te5qEawhPN+aBTF0QvbdqGC60lImdlyK4yWe5UM4bN36h9iHhUHueDVFkaR0ggPjM5iFPlZyWtb
VnNecVGQ2oJENZUZXnDiEpChrJzdWZZtaHDbNgKaOEJtE42YDduArEbnfBPBQVKkitkvJiP+be9a
36wQ9wiGk/qpLzeiu+oxfPY667G1Gl9ZtgTxgszy0nFhZrLNU/tcPmPQii/HxlDxrSYLwjfrS3Xu
m6lVJsbb4oN72eGzfZa9EpKNhJJrwZ75FAhLSTpUXTMxctsDO6G/voTGBl9fqNJzR0MLAIC06/pe
KYISO94a4PFhBigTucC+UZ8IYcUxLN+7LTZEFoScjV7EdPI9rDuR2sH5PP+nilGLbYY/Ky0A0I+V
+psMlrvBwZwbsEos+glo3SkPXlAWfhF+y3XZvNsb/NaFHLuv41OmSEz4HD17Ax6qNbHSDA4BEKIz
NCBkqxNYijNbFwEWx0uAPe1/Af/NZSN0Ego3PTT14xm7ZFZd8Hy8dCqudNpMwkL03qzcgzhsDz6P
GAdkJ732/r5udzHGx29ZvhrATKP+aoEVsuupu+x7ohrEtypx2mNInYL3qlrLxHDXcGuvk1oII/dF
6qKYcM87AbnHXjzCj/pTmnI/WOHMtXt7urbkQviUnOSJp+6/J2Y77Cnv98V0ZCeagsCWWQ5lkgqh
IOKOx1iX3yejj208IpJ4SnuejzhM+Va3MuSuqYdmTJ6RdBdTwkaeO9FjO0G1UG691+5Hs9snGE8L
Qw9nQVKsOQt1mxlSKqu3Wa6PlBzHGXReF6pjdwh4c5zHAfXN0WLjVj3lItUEE0Lnc1q6vnlhraov
T+0EpmNqrnAWqiyc4tbsGVbfSK2g8dF24B8BdCQegHfjAr9mU6uvcfaOFOU6dIAT7LOtQDT4EUDk
3UhmTSI0yEaU+RWS/6OjFLzHlFWRjBJ4CcR36ftiEGYcfe6Bhaq8uMdoiTs5PfbgStxOPCeM41vj
OJ5Mc7pr4gzkHiQVfcY97Z7PyqvFlW3FYqqAjt7CV787aroa28VaGXT+oQ84BTu2VSrAo/WSMOvm
gsxo2/4a2wokjMeuvu5tUKc19yO0s4LK/dUgM9xkIWcuqc4cOtsBSbPskENghpsuZ1ivuHLwPC2i
k1/c9AkgylvhobGtdktfA5WWAaME1z6+hDkXKPI1ys2ktv/Y1NqJ+Iq3217WcC6oakf2GKVJAvgh
nPikrWPZz5nG1tyiZaSMnXB7tDSCNYuw5tSwOhRwJloDqKotR8fVdit++wjqEHuYRresWWyiyAFY
a4fDoKXiASHsjoRfB54q7U9jxcPd6NHZ68nfMcWmcCl5JbXNasmTdW5pbOtavzQ9ghsPs6EHvPsR
O7UVNNW4jShM5AmCu2VJKeWyVPBIqTwdRHydETQze2+60t/mrprXFkAbSkACsoqh1b8DcGGD1sZ2
KcI3wOfl6jDuMnxqbHQPHZYdRP9AeLrc3S2ZUmrlhvgqJS7rA26icNXxX1A40Vv4pHoa+6beNDNg
yooWJek7aO6PlkLXBR9G6I4hJSvv7+JXztqZZGBu0EWo9wfqmjg6YAPlYV86B9ld3Ua+IAcbc9ql
oX+GK/RKY8IsrCP9C+4zimOGdm/XzjlWtmEeQHm02NkzrWoY3PnwMm+aRoXsBk0dkB5oU1tetoo+
iV1wMNJyBnx+/K2XoIe3VeZ95mNoVoPsoBOhvdkCLA+FMkxtjlpQIIBdizJhzISo47BEfhuIt8uO
3BUTNpk+YA4KmiT4Xfw515TtIYUz/4AQMoHed39bB+iZI5CkWWzieowio0kn//Zst/LyBu9Y8ih7
okDofy7lS1+wwlILR1T34dYrlDwXFdXLOgB2lr8GTuh2LwiHw/Qml0u/fFIAqLvnluSWOYnJSY7E
ajhBVwrnkby/2IUNzdlMnMMrPRfoepZ5OVJQwlszU+hNuUION7MiPKvdsf+yfAUViNde5qWIRZFY
L+KY1YX2NguOkDDfVskOlVnXiiyg+24mVY6UN3I5hc/O2Xu8h8fL/Q3K7SAAPOuZPxRaxksjUBBQ
w/oXxPVxckAcm/dv+i+0s1RkZNzCWfb/EQI7GEBeVpc6p9dodYSdUBf0TL314xbcM1g3edlfcNzd
EzzKjm65wmCKN1s8tJsJFUFz8dzQ0s/SoFTyBLSuPxKMJwQzbshLE9fFfFAJfhB9PbL3gLSh2IHq
M4wImOcGcr7tBYsCUVqlsj6uUDw6YUKomgzFCYvVJ5eMSETvUWROkgbX0fts1GZ6m6JSIIJ8uUVh
x5lCdgFsr5m1Pg9SepyTdEWJ2Pf2uJM3U+Q1b4PIW9cTpbfvupC604YvVa6tW66KuGrRu7VZwOXY
Lnl8R778KV4lUjSLxJVXkpXeRUAKdLioRNvy1uDYCnelQloZY9eWlHNMmma3ZSjMl24PgKnGRgj7
gCeGiDBh2zzU2RwKN97716GnZfHGD2bgX4s7xjbVaE1aiY8lJOd7K7UJ3l2k2OY3mVZ9G7jivOzd
dKycmjtLH0Y6EA0UbTdCzBB0SFlBjWcI5QrYTMOtYJIeFW7KfbLJMccc26JRmTKlwviDzivHZcSZ
FOiHIuSY1tfZWyRwyOh2bks7EEL4SPLdNyy1kicVSe3UKqFvuxv7SegU+YxyWbyjEXbmaQ4lgzMm
pADo7Jlxiq4btnCTbf6WacE1UXUjVCrmO8JFRAGpuAZqAOnQv3H/zlboWE8ZfLiIDPvdR9dXqduz
KCVRy+w198JHidbZOgw2rFBYyzATk6ZDyBzIUQSaRGV8k9mQirk3fK2tSjxMbhhXov23qO3xZ9nn
3f7P13hrf8EJclBpgAqN+NgzfLB4g1jsmY2TLQeIbkZXBUZAHXgH/Ua+vlS1RLhD5kaEyzFlqOFr
EwTcEQTdRXWHJT5Pak10yE+Kgo5USVMvnjtkGfOugfSlsagfNWwCUrm7c1SVUGxSF5RZv6IIdAFL
GJ+UYQ2ic64icO9dJPlanckO3jinh8v2Pa/1GWx0G2RWANiUZZEVmJVisJqb4tOzcpNC8a+d3k12
zwd5707i+IqMemHk8rA8mVCc1soVA2p/6kzg8Xcp/44smTCFNrf3z7+9RCKEjZT5OV8EHzJ0W74J
S7NCJ7uQH8QZC11l0XsQc6lYgPZiPcc26+CpwxY+tsw685qV/vxE5aqr+jb4GoRsyNmiwF3owwsY
mAEfuhIIkYfTKdDfSYHCUfNm/IFjB4+9IrW26sx1Jxe4RrCaxOBmGRZWSsy6oB8Co5rczNAY+Yo9
EFwqGHtYeuyd0omQyGhfi9lmrf2OYokenhpQSXL8C4rbpLaegyBDgEAlwpVJFJ2E/wzXJfOThZio
CdxFTpEXrMpbB0QeG+GfFOGZvwu9eCEPFaRGaYei1MRDvu0qtld3lnvNw+kkUyf8WxAvjpGfN6II
G/OMPt/+z/XtqoAWFN/AgFZT5RlTkP8WJ1c63iHu5vypHwpygAvXPpqZ/oZ67qEHnH+4KbJ2rZ3x
MecZHQonI/ZsHuHofn8tQyQFVBBa33t3H4NBMqp5gJ8wDHPzqQe08CLVLVTPpNiYIDv5SmlaZdx/
PnowlhraJbowG7yffhJoDbW59nIEb0nODM0oQ1DOTjntOJo5bTO17TqK4keMWpjygCINfprL3MLA
ldiKyLWlBu/uAvurX8a9CvPRdo6ou63cOdIlX5yjBLNATFoko1O6hHbyLF9ZvKGH4GlHOajPLZ2X
H3usr26hqwvbnZF4tUKnKWgPUxpFTrsK3NZE7qvb6VukPfVTCq46k6hEYxWoMM7E3Py4cpUx9KLQ
rP+g6kYWFyQgMi3Lnq2H/tGcBNvBo6oONmiW47Xa56OnLUc5jy1oCPCvl02NtPvZ3Na9SBOQ+LNp
s132QIP7QA5mhTM7PFWeHl7tyrEPDIqoOx73KfQ6Ky92+8Gb1ux3i+5adTgebWQDjNARf34iPtfv
bLyV1tNGLGJI6lt9gJXLChU5vO35u3+QaAW9UyBoi4QW/xGU41TUiCdeKDo1uZEnnr22xKadA6Ij
O1Gq3V8EIIfIsPviS+zeEUx9YbfQBt3X3pVMWX8scZdQx7oJ4ogP39MSiY8XUFoKQY1bcVaFvrzm
HoSxuPOXvonoGcTpWFSuWa4JuURkj4ip5DdnvEYruo8OMkEi0JP2jOdapFzYZSKEUbmg3wq7T5Lp
htGhiKJDP4zXg6hTuO4hwAH3ZnFd1+4dETiwdK42k5M0ldb/mhKKD7Gv/QBQO1fRdh8k3bOeY9S2
4mLkrTQjmOwe2V6+PAkSr/UVkKv99s3chrrTdAHrMI2b//ntls934bHiuQElZbzvhVtm4M2UFGVS
XU9pYYNvSXfsgEEQpQ1MlTwt1cSBxyk0CTskQjT0vA9O2vvAa5EgV0pMuHDtCf4g21L2s5e7X8X+
+ekgE4QkqYvIxqKuegJxZlAZRKCiEgjfUwT4W19oibqACH4WLOlb1WT/uR8SLnAzdQwXqDfQQSQL
yarRxWfbJ2M+6fMKmhvlhbBTkfhRCBqiDWAehANA9802gZHKu8sFWE7BNgTkGQngTVLWsZSPH/ne
h8fRf2yLyy1si8hzJQKHmdBY4dEcTLS8yNqMKmGHRh1jJW9ARZcspkMRHLHs7mZjXsFH9m/dAZsF
1dtgUx27cBEItOTqk89xOXNDosW1dIMUs9DZvigidIqK8XsFuqSSUpY0vNUthkFGNzQHb7p2G5+8
cyRxc1tNpX7amY8V7/k/qcCK4Ldczysikryi5ja8nD7lYZhtpTxxtxgLctKJTrp4ZweDj5yvHBZM
HD8MjIPCzjOQyMcLVZX0LwCizIoFvuS3uBfms7+HNdsRU8XUlI7g+i5M+/aY44cGKFdGFNnQ5nLU
VnDVrW9Z7fREtpbJJ2sSrmvWJ0rycbWc/pZMah83TVC3AyOlj5NQCPcKdb1QNoSSne2c2M0/SfNx
HOunACJzt/VHaBxSlGJmmPf8R5fiIBt0I0+f4uOL6kyMa39aSMQRaad9enkZlqmaleRaXIlecXwB
65y8pWJupPZfVQJ2MxNFPVVHlFFiBMYPF53PNBFxz+pLoc4p7xWK4BoMQRwdqEWGAaEeaXE1/3zh
iPwXFHx+1JG3hiPenYujxI2ANK6aSgXOdYHBf7XCRAwbiT9fG1RC5OxfIqEXufGlfTMcAalEs8xN
qXRPGhh0qdMWM/9R7RHArlHqCB3aKc2N3gXkusBmpZXhKM7gHxos4+ytpidLy4Z5Pp1lM38MpLDg
68HqrrG1ICSQOWcim1guSyqczXBm45Rp97izoWGkgi4fpUMGlAjcrCiLJVbWN+9jtt/Up3ZZwaqm
6znKKzkZj9GoHyRq8YRzRI0oAT7yETIT1NBaFbcPVPyeSQ2erYtX7bWLhUo1kdknZUchviYXxN1Z
ir17CFILw1LlLZlnxEjVhMHf+iW8aGueWuRMx3KPM7hvgNALFQuvnMcipFUMqGxWpOuvLBviykKc
XJjAFt44adk91Sp9Q4RxL0DRzJQ7ZjTYIDu5yU1i5KR16zZQFPzYFDy4p684uKMM2IP+yEF2bn+b
KbSxIKdqmr3F8clrrYqYYrQnSLsHmtKbBPL7t3n2oPFcOLGe07c7sTByPFk3XaF/XOZFT36Yk1fu
L1XLkJK53JTkTnmcGqyaRBE0nJ0BWXkq99INZLaT1UJStrQisVvvboh/Gup7Z3LFyWVKmAvLSjri
srP4PZHb/kp73r8I8XeZPipZY8Ane8guSj1KtjpptSEYQRpBivKZg5DuP63Egi0sI+EUmjADQxjB
p268Hrq3guYz26g+nymsfpcrZ/0hqdKuciJt6U31luKG38tY8AgGSNGgxoTW+5/m4NSCoQWd8zv4
6rVAEVdFxkLvuWIrWlpoeLvsZCzVeGMD2bdTAgBxMdj7AULUL5VhrqXMgFe/aIhcuRaHlotCw2oJ
H3H5uCW1RRz9nb+/pfYoRfftZQP/6Gi3YFJByxTZLD1VityDGzUc84XXlwgKEh42VbLjgw8674xT
nspGTb/T3ewMkP511BsbgQU4TdkiPJgLarWE4cbZR0xiNSYRTeXwsmv4gG62GXN5a7toMghODwly
0qUyVcyT4krM7sSOqy8YgbN0kV6BsEm9Fg7qzu5bjqATj3LJbYVQARFPa0co+wf7g4F7yJAJL7y1
TfSzQQDlh8kap6wxcO+EAGVTGJhc9LijoeMHiUr0eyH6aSRaQNdRN9bd+fgtBtWOGWiWqRYN/PkN
s7rR/HkEsEQkBNHngyOjSsrp34XPjiL5F3cDPxQjtWkkSh/Q1fMAjKtcgnTjYroJGuOXOCk07fBs
PLPocv9yg9vSiCRktrwIao/LX+YzlXSpVPpkIYZVGUxpzdtkz2FTCy38tD/woPpddgzhrVrtx2l/
iS6Ei0F6hZIEXOc8Jp7qn+upuVh94X2MlZq3EA8eyxUgLa7YfVK3uF1jvvMet1pDZENxksWHd1L4
ZLqeGzYsDor5rjKiy2hanFxVME7LiwTFVwknfdBDTk1G7GY3dFBXM9qdKFVModJauPHj4n0AQ88X
mAz7Djxz0jdDPU7MoneybRacpgUFzaBlQovUMd2ZLIxK+rwbjEfX/5aNaLETQewMbk07RzzXRvYK
JsuWKu+insADAfpPDJR84CuVe6rEhJAzmzDEdZf+xDmwQjhCG3FKaHv43ot4PfXhwpp/CK54vAKW
OvB+/z5yDtHKCXQx7aZ5fk0sqfQmEbBfg7dZD95aiwnGXmQ3C7R3ZU+ApGtcaS7DX1m8T3h9LEaB
6KrEBDiNxj6BgwnAWXMs+E2D5SrWA6wRWaA9/vNg5vqHc1fuxX1lxrAw3get0PsWhThEGW2ZB+hW
Nrd+Wfeg4Ii+iSbZQiqNDJbuRf138IcwTfQ+ht3Fv9zQv0wBJ9SzSEJVYiyAkDHvd+gqV2Z7Mfuh
N+HG7mR3n54EAaDv6aWgHR8asOBDVWpABgygWnXeR3Rz6p9jaiYxJ3vjq9ck+jPBMcmZx8RTRT8N
zfIb2ABDxnP6XQcA1vl35s41q5pUoMQqZNSdu+3gmVCpuoZgy5Ec6JpwckAgehGRTaqUvqD3S0kL
0XiLTGETDopLkVxkFrvluvi4L24v0olGtuFG0nqaSNRpR7hDpU9BAGBhGZGyuwyXra0cicVYtQRi
tHdAh/mBCSIEf/91xB5iPBP+g+iKfnZz2jBIKLpANNL8YPubzD2GjhDiIm6i+7t8p75r+Yrh5qKf
dRbC41LUynMDvOufjfFuDDbfzpQfHfs6oKpuOCRkDXWC4dz3Q5XnoV3isHm5uhV2yZmtEwHjqhtd
vy70HPZomLjrQ+OImwoOw3uc/oVUkAcIF4f3g2JLirOZ7H/KPOWjFg51jtrwbKwOMEl3efT+NCVc
nMoP+MsQ5yF83bEftuznzDp3MNWWKOU00guicG4C6vRmquxeKKhcAp6yUn8LF+5nWV7gfc/xbLhp
yZ/6cUZuQ2BkxMgQhWiHM8peN53jNqtHgN5Vib+BoXnMlwIz+ByptcsViyhV3Q9vskOgpboxPUGc
7O4+cLl9grP9J3i49htsKiEgQ2J1Xv7V0ulzmyOsnqopSaFtBU+AYd0qil0VCGcgnwPYKIbArTIc
+1uSk4JCnuhRQGfxiHpmflnti/khwVvN3sguQGOTVpOI2byIsP4RaVGeE7rTSyA47TeOZAi5u3EF
6G6tTWMQT4dvjc4LizZXVnAd0YRwoN3OS77cC/yuqz8TrJmMSpMynf/LNYmblcYAq9VH+ya6tMEl
B6D1m/r0I++grnbhhY76qiTKau27EhzweLpccsjjFlxhCnM80EVEm8xdP3Hh3Ouxhad5AYP9OKgi
HavCcehl9nyhIMVmkd3GzhvuV0cZmi/tpjUyy8v597PKzhfoMoY1a2Ud8+VPwkyp6xtppdJ/i6nV
Mt0CM509rHdUMR9aBsTv6TKsMHS5fE0xw3Mx4CNfX/zZuE9X1QeXilP2plXT3h4/9U5YbxBxBRMY
zESK1Nc8V6Wst6ioRPBBKXRR7aWovPIWFbiS3pQfV9Bz4PTQLmlWbD+Sov6CWiFiuhSVw0Vb217D
PvFSCZ35c/RKYyHmJrr8sDxnAJ+czgwyiMlFuA83AOyC7YGOpI5qn07+gaF1wNdk7GRH5RG9o6ha
U4cHdwop8eYvnNOSRqxf6rH+cid9F3QzImakixvERagwu74Ovah31kva28fy+S5Nbh3behtZkfUh
YGFQf5SKQv+ORvNf6jEobTfrONb0lohDqptd7Sa9VWH+bfa+Gn984VhNVG7j1UbffQLt9YoFzwH6
zJ1tWhHs3jjFeZ1un1k9Oe9NNuOQ5+5tMTIl1I2vuaPbVG4lR7p0crTRw8y4H5dwZgBNNbG65roP
NamxqZ9HlvTpsseoJ1WK+xcASrkCvA+svamDTaUNAv+kaQ7tWP6fJde8uatklBpbk4xrdSFtHWLW
2SQlHkDbB4BASWql48CbATyg50CERdPZu1jEPViWi3i1mxnxK1lrYkBZuA6eO6xZF/KVVEjrrNiV
Be12TnCTGMf57nlMkRjSuapWl2KgdfO+jz5SNzNaL34jXj445fU8LlofqphBP/sHG9hNGIKRgU1+
oOsipPI7KlYVpLfFzCv1KJZm8f7/JZBLqDawj4ZHcdKXCQUoLPupV2kmHpiZCR4X3ocH+uvTxFya
LwkydujhW51q9dEVrkbqOOZczdczFaG/+jmguf4U2I0BFEJIkn0Lo/CIC9L5Kjr+tPc01yW8Mf87
8VpK23HZBzEPZb7p64WQ5X0Zw2MxJuAYxEdqBuptgUNXi1Oa5IPY0hi3tF598gdcL6sdeZuJ0oAj
yzRGE1ex+i6uro1EtnSptqkvMJbDbhT0UAe0NB4FDM8aEtL23AEarBPxaA++x/3a1CI5VFAAP+hA
Ctnw4kjkPyBGelm8NC935MaWfw8ygIF9RCW5HF9Rbcs9Xk/f4GyLmIXSk//9dfkPMjwonCs9PUrQ
7kOLNGQizo2Wk9bqN413ILJZ0exlCmuWldxreNNohtwT5IXacSGWxKHkHTTia7PAdCNdISc/pj3P
f9O27lGQcA0lW9IXl25e/yONSf4cJ53UAVuWzM5NH0/0zQ7g6Mq1tR1mOIhqd032rf8/RNh4GG8L
ney7n9bw1D9Tkj3/GtTsa7X1fkJFxH5RPIvxYeb/D3HnX1RHCtIPL8IAEzh4QdX342xxp81LdaeC
oe9H1mimV2Cf16JW2QQvlAd+M4W2BWOI65etZDN0bcd1H1pMXDw95WONvWfOMCM6lqNCcymB7wNV
y4Ow0K/AsMh3KwYtd3tyv4sGTCb1tnchIisamV1PMvKzdA8xVkxxCruQKr1hJhaz98zw86Rm+fQE
HKoGUCrnbDW0zG4bYgrJjmKzWqMXuznLRo1SfNbzZpZqgu+Vjvj1rLwomk66/KZV0DPfk1k4i0MT
G1YYTibGdRbkJML+6GRtdusiddDPJQ48uI/PuQBQvTiSIQo0EmuEDvMXbuMFeSogcTNVfudCT1Dz
aWX/dSdlyMOIDGB/HtnziAUJD0igmkQbEVEwWzqgdSGSEk6D3WsVoqUSez3Ld9EmTziZ21+tJBW7
/QZZykIGMH3aAMRFYVz5olqQmhoDCQ67JYqUGgxwG2LI8Dah4OIu2Gq5oLGULhIAXVgzTallz7Lz
afF+uIohMyU7jyoAu9QXOk0YKJbG9QWyhYCRwZm+Kkl5pvZcmu/6EeeO5AzUrpU5uYsrfh3Tq2UG
+p6qZWn/XR7Ve+kpoL43QxY1lBpaaSnLRPCBl4kBc0IxTyejWdZZFYulSFdkqtGeuL3J7VKYK1FI
p2LeonsNHRU53os1y0QHEuwdP/aCpxiguzbaE2eioAOuN1CY1syOrl+4KW0cEhLXeOkdBJRLX/Aa
e+iITdZb1tgFObMVcgO90RAJZ4WeOY1I16lMqgOFieqelXVlu3OPnvW6iedjr/Wn1FTlVav2bHd8
mq2UXKycHdnstU/mdm0AHzLyjKRDUO2rW+NZMdtTFGd+xSqlSEekxJgCW49YLGo0WjTkj/j/1B+z
tFkB6oh23NqFnoHWpw/fNlwyRfppIr4m4hSnclgZmQxwDnHkW4ZBhNSRHJlvDgxv2Oe44pMoI4MW
hylb7GNBiDK/Gpd4ItYrSK6WacBz3fu8nQpqRi6sJxl5HMAlVPVwCE1NvRD0qUY3sImqK+xs88me
5O9XLkXuSRrM/PU4Kb05KEfvYZL0Bn5n3XVWJEBtQH7zR1WBttYBb5dXL42lQu7u7735YYQB+s4d
1ujCbbPujYjxDyaxQClgD6mdhLC+snOebgZbk+Lv0klRVYrrvsBs5EbCpltgl6P8ozEZ6FqkjnMx
XXfV2EuciQ2dPEFTAiroKIRABPTbeOW45/sgVrTQRTb2Zyh6PRg5AxZ1gBooz3D+CTeFvsXXBajF
qAk210qcimO7eZRUFW+CD90MfoWsxVVgPABVPd4gOAHHL44I1ii4FAVe76Vrdidnfs9je4k43ZOV
HNTMWANMiMidefa1qXwFxtecLvkTvvxCK3iD6DlyAQbKdmrZ+6eWuzNoBDOODYi1msHX4V0Jx+JL
xIdLXikwQ8WHq13HuqHwImUfcs/F+6PZuIViTplm+xkHJzQrNCxrK6VOkhbH4puVfh9GtG4T90Kh
MWqlUeyOFgiWl3WyXlawXRk5v0apzRE+tu+zPlwUzOvllT5q04PN0L3ivp2AQwuVmI9n5Hakp2yb
LulvODV9aqoJK/AeBs2VMXjWL15E0PzVzpgCUMn/ghnPrvEQCmtyJMH1xZHZ6fl36cgFZrhMIIIn
zKa8PC7nfQ+fKaz0e01G6QrXlrf2DrXfzTT1fcxc8BWDplSrhp/I2nCMBV74h+tI4jQure2/U/9v
De2TBbZXZaYlB5GJ7CB8rAXaKlxtxQ2J1tyvFv5OLFhIcZqVRu26af7bbWhwKahxPQIat3j8yP2u
f0He11v5NcxBMvFDmobyXXTuGr7aEntUphH/SOrlaKLCnJy6cA42MRiU3zBeZ/GN0qmRoo1Mq8KK
STKUCiWRpQJ1O1vXrJlJyZ4sARoZwUE9SIeSAG1oS1eZzmXnk5nDZ3qlcnxmlFD/kp+JcrCiQze/
4NrvS1vgChEjaL+s8APLtRGhwJWWvNnrP++foW9Bf50Mte0IHHRZtIAJApkNCpqX4GWvl35aYhvY
rkkgOWz6H9Wh9xn4CcYWqpf34QiGCVrojqu8d77cikkZ0Z9dw6GUSVVWEWk7YdbQIG8V0IOW59wX
JLsx+Mv9ul+iR90IHUMeT1xLyTdrrl4zJ1U4pjfErK5UM/sM+kvarq+ZwZYAHj3MBs5Xuk6/WmeN
yORtP4G9eY2ElqNBTME11A2H0yjOMt6EVMprIWpAcSHgN3LDraITCEiXwTmJiZnNG3qMBn9Do6Bc
8B7OSZLnbNVFMoS0c+UBwiZimTjb/H6cc3fvBu8X95suQ294HR3srLlTs/b4gj//Lh4UURSrF4J5
tYW50pM6ueJzir9REhWjkmznZyTliY2InLihsPYgKWW2UPgpfE06DCtNKvzVhmu8niCmOjBhP0fG
+yfyRnJvQKfx3dvjxOuJZ3QkcVG88f8zZ1uCKzWbdR68XIoBQSgait12Q0HS8/1FcjNNxjnnL4ay
9XMDFX8nXTHvHQ01jNeq5HoGFfRizxWInklQre78qtXSHg3TAAHC3OWfV8yZ597W2TXCcpx0N3v4
PyDgS6/I3Eu6qvtEHYGmBymhWDwpFFkPhY9hEMfoAlKYNE6mVBk4OUKLU50ngPwydgS8KXvBObt/
E6nso7H2mQqOIuTE52Xk4gBKDHwITBzJvWxX9MW0qCw86ZxEPa35lli4F3SKWvqU2x/zIoiaKyAj
eHjPeSDGlxDWMvzWufLBms+xqnQCMuuat/POz19A8tquqTrsW5GS41j53H0Yh0BoK+/24p5Ftmvy
CLJ9wWSL8JIH6Uy0gtxZdITuOKM3AB/O3UzlwPfEGd1v0YELEZpuee27AHvx7NYKoUoPKVRfY2OV
zhVb2wvXFuoDgPPvpkbpYa7aat76u50dKswHraWOk70WQBX7FUyGkdXc5yapZiqc3Z5XLJX51LQS
wVqNJE+nRo26V7NwI1NC4ehMbyGuEbF847oM60hzy77RLOPVtRU0HjbObYYW1iWLhHyIrYAHUMIi
Nvs18ASU6EcfEDzrCO8TmEekGMFYcBcJt2dw+E6mjo8ZT5L0FIhPwE8y5WkztcBniuXHffq5QAeZ
LyGGDR34whDQsoXNdSer+v5qHHQAYfCstLoJOIKNEAiEvM0e4rDFW06tUHvLCVl/BsagzSR/Hc1F
rbFgqhWWaznzwYEPBz4BzsJsoDCheWn+Kv6JCyIPWsRnf9vpnAslJT8EuwnULjesby0PrbfEpx4Y
i2PHBVh5lWn57kHW51fRuSi6871UKtptXKk+ngDVj+ET5gmWvHx6/U/h1CpWITfVr5XaczfFp/IU
D3ZRkHynEnWroUU0yQzHchLSYbDzDzQS5D1Jm9FFAoHFbVtIYsUsf+DWdjhnzY8Px/Bm8hINKsPj
UNZFeFZx4esrQwAGFMwkVaCl9eOy0w5xb4FE5xI744Uz9EdMiE4qqk676q05s2ld//LsUxsKqwsd
8hLbwc9GQbSkzLz5wyurpJWQNkrm6MRwGb70fIMJre73idXglwNP/hD4YPVcMzNg1NCJoNwzbzne
/NulABrTraq/x0vMvCandpFAY3Y/HskDfUUFvk0IjBSGbeOD2UDv+2h5+ullLgR1vwIbQP6/M73v
pT1bhNowvPK68jS2qOAQ5QfVbkgSlcn+k8cYoYvFOcZnvAzaz9FUOvMp5hxaOtM6WLEog+iLphSf
tfPLrlULegId/PjjfOm2rch8E4jQD1MpFbxM7jfl53IXOatMdzBtZoVwpeBdXU8G22jn9Wv9g5wr
0arikBhrkdOWMaKQ2TEdraPX4mq/0T/alvVm5O4tkfUyCKmqk/NLKd8n+PfyMtqiF+kSNgiFcHzN
aCkhH0LVwvFDp3Sn85Q1P6o/6fwTAvMNeltZ++P3idLFBbOwaklQkRR8x2+bJUWfBPs7OoTNH2Qq
Mq9SePTEOzpYcH4wPVBL2SeWoPohlowVuzTteLSHdzsTLuaH88RCzzTPW1wfTD5KzbE794oxiwaP
RSP0Z6+Yw7ScstaWznwRnADLaW5koxq9OMCGz6icUD+PnqpXFA6nOBeZihlASOZ93AyzV7yf3tLa
Fz77FmQCujOTHT8pw+3e0UrT+hpJLn2wpn9nmNoH2QhGS6hHyVstzCqDDINaeQYi1hImfuW5Wkir
9ldnEzTCXqrOMaUb2fFkSUHzMvpqA/34AgUVFRmv+YrPbdkuCKw+b/BmEbKMFyFLyO1ngkObJZBx
B/XqVE2Ze+QnpV3rWCMuOP7eQBZYdutqhAw+fjTULJO6fJnpnGg2QL2DEfvCxJszv15RTXcz5YBZ
14OwyW8w/ZDxcUQQtCLpMjNxhi3V8D/sFf/rK5neKPDW40PzxpIxrgaiwsKU1z0CAQvcMaxyzmoi
7B0aGfRHLmXvhMz1jBiX26mzlq0EZx5OvkN8fr40dFV5Jbm8d6SQQg+0lWZAHrJzDHVQ1GpOMj/n
Qz28ydsQPnVfFgZryY7X6okAoxS39No3QJFzGvusCIDihkWp7QyxoOJX+NNb4ZWukdaTGuwQfIoj
LB/e1t8Wdep+kYKmR26plxwhqJ75mAyK8PXEJSBLN+EvjGbVKNzh6AV8sp26Tz8Hp3QMxu9rS4Nv
SveFq86oqgGpsjOgd6IP3SaKwTi+7H20aRqb+hQKU7Vy3F16gPZIq0GtpYAkukTiLN6ql4dZ/KGR
orOFUxgA6waEvkcYDV5R04kWlerYzqh7b8F0bu2bxlmJOqt/gV1Gh6SS7UmVpTlD4PcF0+Ok1KzQ
DQ3sKcM0wpl1qowxlenOxTZkoj/7sXLj0B40kN0MgryqgCHgujFc5oR6Momw/Cmbpy9bq+sLPc4k
EjMai2IIW3h7z4tQ9jbWj5crdLPzie4es8xfDSvNo7Y9Dg8KGDeSntxDwAb38LhdAv8vbBp0U+lz
lZyS/wY4Nzm0BT4qusyo4YYDU5Xb1hVXRTo6Y3EDy3qKBhY2iwyd9msrjOMPKEceH8Dc8VfBx7Cc
Craenr2NfEonla+NRys8IAnVDp/MRL57HamZ2Rrt9Cqp0yjxvVCA3leFonG9L9cxBr/D3Wfj+mi9
Nf65sX51kPqyh96vZcSRmc5TkbqgnOCQxWGl0QGs2TQfFc3DmKUc3VqBsbmFQhgpSp56v4JjZqeo
bpFf4vn7OQxs1n5lDrgrXemoqJ7+7AOhFJOESoZKUr1s9OkZzmnHGXGFzW+2H+z8c2O1qTpk7oRt
kW1fw2TdNSwFo3gu+pAR2CTtW1PDwTC5LNVlucsKs6ftLdQLRZ60ZqqGoF5aV9wpxExG5jGHPiIS
c8io01Y/JhFO402IP08w8Lp4rzhkc5HrFv3KkWDdhVWpC1cXLMZNQsRL4/BstNirR4fbooFHDmGz
XITwYJiCphUYMbRXC3MlBkZzJwkvEGYzAHRqGzm79Z5nDFSTJtdTNxk+P+foQZM2ypnGR6BsWf3m
bt0L0paYev5s5uFYI8D85TFXdn7PEdeaCX62J7BbOcjUJlVGpmZzcWQn/nUn3PWfkAlViV66vTKl
wlis45/kCLBILbmT/R0FMQJPiw33mq5LuF0lU5DZdjiM5K0jdS3oWRzsHrTOtxyZu5TCvJ+dD8Yo
tf3FEeY3kN6JVGKH7gYrj3rdgctH4g2NuflKE2Pk9t4AK4SnfPajyAWdlGsvid2o51lfjSWnrXLe
JKeIFcOgq+dN2B9+9tGNIobbq2E1QK8S7jBjIkukGwJORkhQ6nJL2BLVKIVAF4PPNAmebJZaKakh
ZMXf7lhls5VzmSKd7i4oqofY+rjbCUgRf0MLyuHTmgfdEXw2YhRGRdjtdnTqogfuKEC6hDqM0DU8
VNR2zeHiLjJU4h4lmGWGDsMF+YWs7HVcYjH84x8hzPAjNhZooLG3cJz+aifCOK0Yo6Y6ehKt+jCX
t6guaaSzEiL7IvHMwNokvMfhMLHRxWIyH/jmODbgStJV1OerBRhqJyb83PGpNRI7/4dY8gY7SSGL
Aw327LK3TX0OJ3d5y4NdeJ8QsXZ+njmmJoFiwVmMSrYGcskF5UN8zRGS803ZjhY0oWpKMYdVjWIa
ddkfNe/yt+vHjjbpjm8KCvgV+yWix6QId20J/lWrZ+uJg9NC9puX20LDfpH5cUdxr8WRb1CNUWLX
Ula2mY62aK/1vy2oMOEBUwk/QsaGok+tvLfo7YG3ThvdSm03Hjht916McOM71Q7lPSmIlY+/sFP2
+oS6bCHYjmyR4RLpk14zI8CoGkcmFGa+bqZm8QmgpKtLQjBxLCAuRi0xL1TTrXKQqPEJEo+gWRql
rIpnadPGweU65K2O5reS7fkpjkJ5XT3m/rr2SAG5u7VVwUd1I9r1/2sL8XUMA9g++64t7ftoZ4nv
39F9z+ALoGKc9EPbu8YyHp4KIpGUWww/hxYuy751AoT6of8Xk5Fvg2X3lI4V1QS8fYZd4IPJT4qS
cZ/Tz7NhodBM5gVV2QQu1z+Aik/Q8/YxKrgZoPV3XwfoTzZzwa//RXljTMu7OHgWT68QdWISxdFl
9A2wBRPacAHlZPZhQkeGO6yD3rXnFLgXzMrOjKm8/Y9hE3uyb1sb29OMv/2MHkGBFu6HIZU6r/iW
QfMe6zHkoRWZATxagr5rvhkccnSwtdzigNrQdyjMUjbobxEyx2thYH8DmfCME3i0b2R5gBiC5ezQ
b7cd85P9XJyzRZZRi554yQiRcxw1nABkvRQD1PeTaocLUPXlL/+FK3vf0YIwamyov4/oVm2ckIe8
Ih4mvtwjee5dT/U9kYI4K0F1JAScAWiohIezHQZLJ9l5/5iY0Ivq9SSnPlMzpFV7YD2SAxFYOTgE
v35EEmUUlxbfBkgVr6uApvdiJZg2x8k0dRpwAi6deWPEHG1mE8P85Uk0VnGDYb8SSj3m6MqWj2jt
1q+66PRj6AEUt69fGDuC7zWa+LDSaayBC+lxwtemoiyp7vxEGxsHHSEulpKB5cll3E00/FETWAsB
+NMfYdPdA0d7YWsYt0NdtNRDWEsSDN9USPpKsWUSRFmHBtCj27hfrAWsshff0v0XveK5FWr9LYcw
wD+ikTYjsMlPgGjUEzZmnNnTwqPFnYdG43GaIGzo+mYn+7Uf7y/OS4l3Ygw/smsMTneKGK/tnw4M
cESKZkBXqhDmcTjj346d5P8HM2MmJjwaYFa3/zv4p383FIYhTPeyMpGRTiQ7PwS1cN/Zx3ah7GR3
IHihVGW+jyT5GhceRPqDijRrrHofdrEgNYqZeZBpg04up8qBckHtFR9kffyad5f22jAlTW2e/2ef
hIXlAZz3PCIfK1KN2ON5F2Q+H1y/6ss2tudhYMocT7ckxZ71NC0DxGpq5p/LSW/ogH4Ks1L544Kd
0f0Bkv8Fk5y+2K1oNZmsrVB4nx7SssjsT/rM/IkjZjtym3oEmr9wyTX9OY8xPtYPBlT5MeUUP1KX
OKeP0d39DXCZQsupbb26ZiA3bYjvK9hN8uPfSN7GnOD3dOmH3+6KDjD+jocdskT85ASWPXJeG6lZ
ieLZb9nrxm960Wyq2FX6/Gv0xsw6sRAnjdkqMz9emL+gczX7GRCm0gOHFYo78UUELqa2C9JRcuKz
R4OmkHTP5MWVvlJAuZOjw2SxqHjPVkioiysHWtP9vehnW6jMexfOvldmSwlPpBOi58sauWKGAAiq
qUdco2q+/8/hZzZAvW9RGa9N5E2kdYxrhV0xZRPqRAsTgG6OdFqe40hNS83KdRMVem9O/5SzieUA
3n5/dpgq5Pwnb10HohA6kXL4HsgzUm2up6z42W+6s0u1MNbA3Et7fOMyoutep1u16iv3+lg3zxxr
V3bxZiwD6g7n4/68ktsbWJp30heO81EfD+VwWOLeP67alg8vchvV/6WZZxLjHjvy0V4xDCmlgsPt
82k0lOvbAjb9uiHOpkSWielPScyq9IAH3ljJPJApq2t6zLI80y3TD4rw17Wo2a4+XIAdmeGbj/rP
GXNcSygemZbnhVYGFbZbvu4eC81C6k71bM7DLue2DtOsR3uAfedWCgPUnnSpOeYAL+BydVL7zLb9
zTHD/x4nHpBni7QNimG26N/1iOGNpH/pQ/w3z8GcAemIHcEdStA+3Mb/pDtfGVHezk+D5avBaOwI
JPh+bHT0jHc9a/fDtEIn9UkB+fVZbMbZjqIGc9Ds3vVFduxkfdWngjULcx6WpnKPhmtEOb37b66l
lkKoRjUJtQoTlbZegnjVPUzNd2N9j19tnAjzW28HtkjejhXCbhuZeJwrQ0Htrk2uhLKW6JNWaMEf
GsHLmg3bEKbHIbIZJ8LHNzWvBWJ8ZGtwkX0bpxGTqPiIwHyXWe+jfdyWpvIb/ThjyJoAN7zgl+Ue
B8RkgKW7hXnfuOXjhtzgzLFAZ1m6Gamp9CAfd/XlbiVzXOklLnwrUfX6RujfAaqZYxf4PN7GebPL
2w/bQNklWn6N8LUbGGoE05ndV04w9xG3VeIzC9DsCMJHzemL6qc3/Rlo1NJ+ixmWw8nY9o063z85
B1DVILRMfvDFb57MbZ4Y5jzLzt7OIuxwhcNNtsgz0YZr2Z9M8NQcvW7OlMYj6xd4survShLi4sO8
DwOsgncNX9hM2RFquBJ8mKxSsLrZEdCgCnzyNoyNSgPr2/MHLFbyafVroLhLbFh06Uf/yAhDeY6y
hT7jecCRFkkudJ28a4yAASCGk/0OpcPpXAM0cIaLC9p0dPGLRDh12twgeQyTS6c4tNzoN9SJfrIP
b0gGT+9rQxUM2HVyz+L3nwwZLGxyx7w12wH9EoiAEiCzfHaX/4LuuioDGdSSXIuT9WjYnjV3XHS0
T1la/ykMiir+Ok2niKH/W608CIMgCFbavjHc5tgEGZ6RT/Egu5520vDRfxlalUAjblINA58jDmgg
3h+gItQ+mF/WSka7zHZFJ5SmAxLTVFfgENOd5y21TcIdLSbYrE3G34k1RLhAqQmRst+Keu+YLPlc
I9XyuDJRIT7k6vzaWjYj5FRm5VydAToF62XnPk9k7w98VfoJ0kGFRA5GnvRIsPXj+aOAT0mqdcK0
Uro76KNOFlLSH0OzN/aMHt0dUHk4SgwFkM/VB+XQDGz0yw4T7ZPdDZUC8NuMpgJNC4SdxFE6A4On
uwhDpoNBzYatuQe7VIhP5tYkALE1GOVhMsz7a7RcBd8PS0xyGb/rGUZBZ1IVP4qAhmOE26zT7n6V
hxggYaKy/zimhLmoBxc668gEmz0Oi4X62B55qmo0RdCJ9JZiBkSrHMrZz+54ZbP3ZxVZnjSBQ44u
SY8o9FtOJdFOznT2bA/qKNmOgLeSvUlaNlVVnj3QykWh630o5HKXICtVvtJZZd4AhdxOCl4wrp3m
W5KIb4/4XvLOWjyOaQMfxwZzOY6ewB2LSx2v7YgXj59lSw3P0MlEfXh8vmguSVdn2NlgzQYUGo5/
TE5u8UK8l79PrKqQIwy6ZqhjyAvs7VbgD4hg2Ymq7ONCaLy5eEfUV67Odp5QImY35MBlgO8ISEJk
zV8hKjZ2jWS32yuUgie7w7FR2LH3pVsilmISWGGVpqYK0A0lN8gSyCIGafrUwWDSke9u1ROO3Deh
Kfxgfvuxz5qBFj6SCNyXWbfzjo73tvYQVX27tscikRPI1HkPbNbfEwULNocrBTsV0qFzXVt/G5Ce
WEpIs26KLgckOlBVZQNlj0ENY8DBtW/0mfSBxYfwA8jEpcg0OXluyfyM3H4BkgXDQ2N6Cc1GGE5J
IoBBQJcaPgzMbTN+/lMj4AUsHG5saHIrpVRUmlpU2XC2pUCwYecTrkg1Q3cqo8e2VQtUN6B9NTlg
1pUyKM6ubv7NeoctA4Sen7BTObSY0lssixxVwIK4Z6SD6qDI1/ktOrySt03l2vy9+8L/TY1e+FZW
HCQEPwJhNy1fauLnhDY9HKDYzzHzUU+SY1Qa6iih8kivLPHyK4Sj13hLXWOM1itNkd+6kPuez4kl
N5IehHLFSnDMpzIq5NXKc7fiamRIfwFlm6WILaUYwvKtcSI4xPV4P3sMgzWcal0aqjfoRcwRVmxk
baZg8jJLaZGjp7MZsvYI5dZlkTpge+PGcNDZQ7SKWbG09SXYnYWf0syUuqUlFGNp9jbxsPfd6IUT
CSNZAh4DiQW7fX1h+PQBi8KGb9ing/T41KWHlGZGFG+c9y0TqztdYKhiVpn7kbrgAuVbrkhO+9h/
FcVLGq3SAcPgp7z10nvGtUiuZ/Z3+kKAqQOD3+dkM/I+TIKkH5asgupcxwnp7oMagUhIGXmpOhoJ
gLEnccw6D1ge78qArja972z3cxXGrzFBsYaeIPX9iHsvFIf51PN/n7Z1AZ9UKpVQS4Oly3UPpKyq
RpDra5M9t8rl2t/6su8Ak0iU1CDzUcxwXAUSBqOi8tM3u0zSpmVCrYRpFnb6BjSaqayF9oIuuejP
83yLw/xp2kA3raRLRMsEquqvW/c4zAcdEv3nMramHftFA9mr/RiildRcFb2pXPDQMInCNFAN3IPE
ZVv8a1EXsDeT2EAAp5PjA5/o8GPo8EXEqnQdgR4LKvJMCJTXew6brhaTUlKf/JYUnFo3q8pGanDt
Tr5YZmXvL2HxSBSPaab0sRYwQGeGpE880r94vsVE7XDoZbUgntzeTU28zk1v7ftpUR56m5O1oEss
GwlRYQy3a/dbfosniNmsQYO9d8E1mJImzJfGbPeNCtH4kOkuYHbRNsl9t55hOPiHm8rjruPYI8vs
/V6fbdlsq+1nnz0gzvBe/4AIJoZ6o2+NbtwG6QVYajlMab7mHUDZY7j43u31aUYnH4SkdAPcBRI5
03FcaXSfFcrCwC/WI2EyKoPNfU2sTspHS5XoU+S9euoe1MzwOKLXvqaQFp115zCoBOOiMZLYYDC0
U4rg0wGO6mwC05Rqf+xwpxa3lktVQedSR/+uMFjCpfZy3bQ2CtTtRcJKRogNKL0TCHri1ZQeep1z
eeyNNmsu58uZ8//hMLrYjc4x4uFYUUMDBMlj3Kd2O54ozqiGAa5YFA19Pa7h8w+x/FevlYijTvoR
7VBiBK6kdoYsby+4dPOfXoFbioK5EO+efRrRSbS2+fP1u45DXsAI4GQ4NEAE16IOenusxBdXvKBk
zneI7w6Qt3PrPDXTLUXo36O8HIHJpqqJGeb/lX02iNEOqNc9uGvyZzEZU/Vk9hoho7bIu4KBkWM/
OGyToRH4rry6mNri0PnGHi64xV8/o1Otd3v9HGgdQsDshbNsbxdC87hFV2C7RNG6kV+uRsOIHZYA
5ba48XMsFlZOJATtn2DOMFtRSvXgmOMEYAWbekaBypWQXbqcl29NvMgrqAF9h3NUGmJEE09ATSNC
/b8aEgKopZcfOJhAXmqTdtaN+13peC9Uw3Wv8UeSb40yqqExFkF6TGoitfz4VZ7+AS5a0kfE9GGv
1tCYVWZxcJBhH3kJVJkwVz8OLh7FCXBEPoxNDW40bIVYMIxRXDEGmyQXE0b4eVo+S1yF8S/5gx1g
LxNIvlpmZRJxsgCcAnq9D+j6aicXEKqG5VVKe+3kkjU/KY0Oc7xPYV3sZRAWT8M4bmsT3YiPqamA
fOJOjRrdIoMnGFzRjkg855q3kq0M5bdKpePXCC3NFYAdqLOYaHcbF51aeN9mOdAO92bouxphnllL
ufXw9wvG/XOK2fBxsQoc4Xy8RE4bWTggb6dHT6lcdcFUrX/ZtBEc+QM4GGes4MDH/XTL8ivTd3b0
e3IVtKveXUOzeMJ7RFkcb/agzNSBvB0ylrKkz6XM6yXbo/Zs53HIReHYJZv8eYgC5HFMNayXb5fX
WY/z+6PkGbKtrDyI8GXiJn5Bc4TOCzQKTPCaQBn1WXKBvGO4PtCE7ZWAzIaevs2F/TVYAtPbktNO
5Ml1MJ2Crn+SQoLNk80mwG3T9h+deEuKwr4qzikAH8upsqbDX46dAFqWDj/5HTLBqKxMrg6HatZ2
pucZWQQ4vGiio1+TnIcVWjOSbZPliB8ea98SJear+GEJjHhCcxtRzRFeCRKYttZdk1kmxnrrrc+u
2dZYWzhFhwdFw6seohM3BweFnzQBMqcnA0Euu9fT3oTNvnGrhkJ1MvqZ+zJMkcnLk/uWLrluYImJ
qBCWbZeE08ACL/oD4/YwkVKnTd2LVQ/qZ2/rerrPlcetnuTjED9jsBpPXr13AMZNBndpK4fZQyYX
Q/APl8dJUhDH4EfUu02q7P2bpkqqAgYxwNlyGsoljPBx4ANVs9d1YKTwsKQvNSIkRPcy215eypyC
N0ufJ4zE3sLHoU7+JjDS2oUIXq+9TF/b+Cv1VSWpB/szI6WYGWiYJPog906wqzFm/n3v7Qk/Xv75
YxYAYHcuO2NY/IprMrTYJfbeZJzys2hBZAjh2Qb/uyxBiY8zxXyCTaNhOTQ+TcfD5iuYU5fLhm5P
ljAsVTsxTnrCJric0M9p67k8Pj+iF2UhJbbl+KL+LE5rb0J1ujtdsaj3sX0XTE2VWS1rN4FZIxgg
DmlJj+nhjc17FNQpzJaeIG6iBfhc0uIg2H1BuJo6G7D3bx6wE7CsR76efNi6vAmQmPPbJP2tj8CQ
qTkZ0tIa+J9PjGcKq7DLsPP7LWVYMv62CXKmFNMHqxzG/grCCSF2qWlMAZeNegVX6GDxO/Yx9eiT
t+CL/cpOMZrB5Q5o31fai6dWtCC1Wnw1Y62RtZp19Ort23amsX7uorOa9gxFlTidF0Cfig7yRdmO
w08o+OT2ANjXjMfctyKBsA5VkoWFrLfcHHk/3jCEIhuzFACaHZ4BDtlfs5Eat8yGKf2rn04SyBTg
U3vwXCCnPU+vtVNfwn1K9SSP1rOHfSmNwunjJ0BcYSr6po6YlfORKtXMfn7k957TeKi7rvO1H95A
QuBo2ntUSX8sTt17vFGsbS1OdTTtuwuaVwdVo7iKcC+rWT4XmShmrjBMma6dZjINWZmkEgW6atIf
Yv8T92mTOD//xK9MdC5BuyW+pa1mQm7O25ORVGx8ZTdkDOReKYXZyAH8BQTVsegHwf3BoktO/GWh
0+KtmmhYGQh90fE2ivYFgkIFVQ7QdMQk8BTmIQV6D63coz1A9f9zTGw2ht5MHuf8Iu/xamHglXN9
dzOoollNAiFtSQFDSuXP21Dddw8m+/vC9DtKs24lxNFLStO0afPxf+RCpTp4luTUF9bmhANUtWaO
9qUIMnMFjnCVKSwz6pwT/YFAKclAT2S9JhhpkKAyfPaKDiN/mRHmoYUBilW0OIaExWWiZ6vpSh/m
9KjESFa3N/+08WNVwcXz30CFtU6KTE65pXvg23XucFG21HfQuvnOreeHa8L6YcEubCaJJT3efXqA
Sq5BfN2K9iPCOzEthzGANptO5xmPXhT0dp8cQx5Pm/sEeA1dZZ282nLYg2h0SmgOjAqz5cz6uUR0
1RiKtcK2MYXIQi+A1s/EtkgphGaPsLBQTMMrS4Ww2BN2XX2Uxx4pC5LJ6nxmgjekTH1/ezpzgusI
L2/vxrfbkqMsxeK3/QOxCnlmtHX2oGKVqwYG0HlK48owC8j8+N6ylp3I1qxWsxQUtTIngEm5PsMr
uaqZ6/Vqhd6YCm395jeaxIyrp0nDgV6ywCQaFW1X4eug4nfCU+MxcqY6sRKyY7ZNdpHip0Gm+vCT
/Q7ZL2uqcKih91YOKkPFN/JkjHSqrc6RAN/Te5SPPnVa699Nj+1Gr/s+xX0532elk1Vb8wKofeix
bPVCmKGGGxnZdBsBY2fbc4q3Y3A/xzW/C4FQytRGcJZvcsMGMmUk38Cuia6SGuo/p2v1M+RIGUm5
71J4+qg7vmwK2rSct5Nlu37rlYuVMDYes56vDIrIHDh9TSp6x4EAS4KrzobDMJeBNKbdyKGqq9Is
B1jE5uVAQGmvV/9RXTEz5ROWKiafQs8NgbGHTJ2p9f7U1g12d/PlbnmiP3QmFGHWmHSwgRRU6CP9
1ygK3b89Ykb9oiGo0FVt14/vmZ7jqIzZ73FZqHYZzluJXhyeJO0TT4VvjEWOjaCAD6K2FYeAl4xB
AwWKILiehjb8M/j34MX/UOIo5QrYPgC/5c0kMtaVobs7B5eUNxQ84MR1jyMwIUPxFn6VTO7Pi97Y
TqgU8lM84w2U6mqlQ6U8yyDC/v+wthYvlYumhHbW85KeDRujlFDapGxL/GUUkUg70bU6G8qmziZF
PfvEBelUu6c/kuSRbe9SAMrBVxkrCvsk5jF6IZBIMMsanKHbf4LjpZ4nqIMWUg9MkFup32/wQq8d
QkcFll35X6Ts/GaXTghusDOsttqMCs5Cxo1b3tv4qbfbdai3ZV94iCDnqNOPhLO5szbOixclyuPE
vBAcTPjC2cXxa69vDPA+YfJpfuizcMhpOqOOMAQVCZ9TqmY/gM4qEi435H97Cla0F1jyUsUjw7z7
UfBVdyoN5OTgzrd7cuMmmvYAUDYySjnYI7LHH8jXnW8po2d3Q0Tv3bueJVg9rJe73zudxJqrGsRF
Z4MvNWeVw2MhPxZv/r6kBYjQqDbNO+S+95KejOdPLs0wFKHlVHiamuyzfFWlcNbqjzHKnfpCoHpH
lEPQKuL+fadYh1LwMjG9dIGZ8rzyTgx2Vt/Awen8LlAk79Sb+d9UrzGJ2/+uwk6Ck2BQ3E12vFjX
uwvlxzmxTYP4mn5xZtXolMkCWppi1Kbvx3wgXb2j9BnG6MAElYVWFdvviS3i5xImqn6pzAvpzs/5
L44+MePZ5YEkGQCXxI8xozwEk20lJj9I/ELeT2zM01CSv4LVlVnEvsinVVN7yJm5gTRFV4M8jM6J
dQTdFi8+bFUGtmkFFzOdVgdqtzYjV3IdPPXmOHttYcekPrOp8AkWYPS2PPT3vK7Uy18qQJjxgQkV
wBnqdP94WfaN3DngjKeKhZgc1U8xVtgKEpXAZv2ndxJ79j6fZmht6ozMdAMvwVESUaS9STE/ViJU
4olJZ1ApB+DO77+cBfCkTjLdI+g9extKajq9ObuJEuCsXyRXZn11jqMF7uzuE5mnxu9ruXo1ZIT8
3C09skdRXFHPni6EdRyWQOgED0W7emb0CyLeWDZIEM66/g243xkxmVAovK/1aTM6ISWxojhQ9/1R
y4N1F/NW6RJkffSZLOdo2fkMr2z28pnLPpkEK3xK7Ntak4EwCKH3G4IUJPIeOgzivlq1HWKs1PUE
2Nokvmfw52d2xwdBjiKA2Sh+rvk0x9FWGmEtjiIsPQwh+P8kKpvG8sHMOjsF9TD+oW/q5i6o3f+Z
ctAYYAe+6t3zcm4KMSvDtUoVnxr1oRbKb1SH7hrw9WFANo06FXoe5CZtty2wZkRFyAgomcuYzBZj
7yz/L3DcGxVKlZ0zwEmmewm0VdpgpnyK1JMeK1NaEdBHb+/saiz+oWA4//147jDKZ9ZoP5bEttod
J4T2xFua7hy9bR7izhx8Ma8mj/4sy2QjNKygZ5pww721j8QNFSInDPouSOlKpQpmwciBAtWj2Tl5
fKUfX9moBddwr1gBKupjeki0MYpM3O/MdhwpSjvuX9oEmG+U8LuWEQQSwredBD7mJTh5NHmvanmQ
YsoLPFROcu7l91cVSek5CXkVJkezKZu96piFYQVkkdASRyAGDiJvSI3oTLSZVkPkZwyYg3XTksQe
KF2h5CNRKDkSSQ1vUwCxTI8z1Rn69jbxBBTvxKcSfSWvkAAeV9zNprAhbNuplXsFUeWqTN/8ZmyE
zeXF5rf16GHq8V9Fe7XArTNKfwEq2cnbR0gQFiK/7z0BPPMax0fnrpKPH41gweK5QoAo75xezOPt
DiBSEY5RnZwAU40w0t3etPQQizCYnbM2rDiML8CR1U1JWY59eyQ49vreqdUtbcaK2hI0wgOoOKZX
XlVI9CpWexdwzfNHrIMNPWxG45/AU3yfGPYhmnhLb6cUaefHAAnOTQ5re+J0EnCpTHN2TudqIqDQ
MCxWJ0hyATtNlHCkXpHf91PrHIJZatXn1risQdcASkXEEJoVyjzghIOQfG2+9iCefmgUVfTSgwJO
VKUvtVv1e1Ju/MDEVupqlgWc0CVdx0Y7Fj2hOjiwigLjsZOmvgVpBpjmtH9Qw/QKYeIjJQdDB5BL
nWtV1GPpPzDc2eUpDYcaeDImRK8uS6Ux3XX5/BqvCYiMi6FYQrnU+uqSbK8N0vvcQRUuM81e4eu1
OtcEESx1QNExxEAj2Itj5bIBomaxE8w+wcQRVlswlqGC4DLZLqOTWoGGg9gM8ORJ20xP6bHm6g5C
D3CXYr4wIjQ29Ct2MUEJd9bsflAVUgZ8m2gXbk9ICQhuH453cxCufKPA4lmRFAQGKhfXg0blQZ6M
rft9dK8LjeUEBTs92E8KTvVhv/Y9L4sJl2NecnisBywEU7jmQ72KQuu8XJlNQS0L99B60FaXw+/2
C1w+HBRA0WYKpsPCLHqiLQYkaruGPpvuU4xffBOPmakD4GHUKzf1FjBUdd8/gNvpDcm6wcW6OVz+
scGTSfX9souV+obIjuY0Yla7ODkDRKjia8fvdsconNqJkSvrbTqKVnAXrxgF4ptxZOAz+ox/Luvp
ZFWIB4pm8iH+lpJFYkJxarZjuiMQx2V+P+BBaWOEwx7jbtO9BJen1pK5y8G+1O0f4kfWhQw+Pe5E
7KGoJCHYPumzQYk8pd2XgBPMjcGXvfH09ELdRbuGfDkazj0LcwI+Fq8kh5bmSJCOrM570UGyDzlH
pjvayNJMqSK4ckFPhRAC5aEfoB9h91U8lUhmex/iNMLvXLjKHx0kz+nQ38ZeebvhbEzGH3CvSsX/
Frx4vsbG5iLqtHLxVh9KlBEJ+PuwkX6OZ92XStuEQHWuigDJcJ40coqYT+6s2AWdHTWy8LE6dAzt
VbxlMFpEHQsCO1M3fh/XAd+LXDBuknQ7/EUMcJhEgzaG9RKlzDVpnF6swhRC+Rp+3Jg3YBMt4C8S
hOwzAlJPVyZ6mrlDLEHRDM72VY6qTvh7GMOJYmrEAP4oYhAzv6lLG/t8oFJHniqswBIrDeovUWEB
r3CWUXygKSXEkPHyWC/zpuCt1DvCh1Hrzs7hstFzVBfJ2lfsbnaTKUFtpKalTbq4ShhELKgZysH1
+r6dibRPeceY5fpQfKF1ac/cVChUyRzDwUGk8nyFqfBYZWKBIJgpBOARfmKsc4sP8rEoQLFu5Trv
wBuYKsNN/ODIbx9DU1sCOj7sO69DPi9OaRLcDiVgm7xmHUa237zyOAypacne9Bdk7eDlCySGYQVp
bg2rorSDAq8sMADR4LUX+4LB4kzIbm4zeoHfwTfQpcrxs5mJE71jR3dyYk9RR9FJ4QFElzZa03aY
EdJ28BIhyOogWkxxZ/4RRpU7GMrEx/jmIbxVkgJAJ2C9JPRQRYeXejFhUnv+08gFdXer0rqZ/F6c
EjBbg8t2aubSa1RYee1xSrqsmzcf/53v4nENRYNbAJWKmEccDTc3W+6P+sPPjcUBmj/EQFMKNE0B
gcnCGESoQcu33rWSo1LHkML82YEahjYU7R5ir0FWkJOc7239WjKMr45BHMFx5Bxuf8Vh8oZUkHqw
c+crAbVcc97l7SrFtmRR8X0sqeRAQ/L390GFDZxU/sGb7MbT0oGzXoC8Cf8c+st/pbBrFjDihcyB
ZbeWYtpsBrOUhp7ezJyKsPRJGVXqXsYAf4i5f1kGQ83IcbEUB6Y01cnCZnteLumB9LbHPTdc5Qbb
P4//5wrhtJyBD46jmvGr8ZLg0t33C5SC2IqDO2jtrJ+HbzvtaB0NqJB2n8EmK3jtCXiJ9VLbrVYy
ILMVHthM9ZjbEmCx4xknN0C+2X3iawyP9SPXYPe1EcqG0XdSboj2Sx90YDAXwwW9SiYqUwas3jDc
UDssNZ2XdIdG+7zQsUXKOl64pGHisPa72zjuXz2Zqglm1AxQTqMAXuUo8WmCcG3pao39nclPtQsh
vvS8PAIEHw8sUFGPiJFFwm3XOlDrhotpeHcSZoMZ14vreaBztlySDd8rTgzL3+t5ae0GPtlQddjq
fmPvDrPxwfia4/rxyyt6+2JYVVxjzwe0iwWC+6innogHQBmZme6NLAq+k+rMUwYdXvIqJHHPJ1kc
KcFO2vUqSDcEbUc8J9VHvSivVAP55FyTWu2/9LXGvRU+8k/oiffARi4UNkHApzXLQ0Bo11weoei6
aGPnVprK+7Kiwh+UcSaOC8PgtEQf9rXoq2Oi4yQC3+VCqE8TRfKqk0MqFkRmBhNuLxTlLcxgETWX
mK/bWnax06q3/VgMODPE3Lg/Ry+QqvcfgQ5lNUiHV2uG66S+Xlq1aRuh7kSTH9xvAAkNi+8/0bzO
XnI8U5mvGJRpwSftzmKfgS6EtD0UZGnhQWJS75+zoo03NIOK1IlvVykibHybGNkG71IxJ2RtylWt
DGrKI5knJOACGH692z0dqLlRR3/lGEbLxhpBsxcCObB4+RLRyQNkiUW/hwkxMAvmkcgOUBYsPX/z
J7bVR805pWRk3mpWGS5QN+qf8Vd2TXmmIhC3pL/7j5cR/RM+ko7ockavfKDHrkDd6OEixmTMmstI
BUlMN9AoQPE4o5Qs9DLG9sPtlLoODLhLhYzYcLVr5Lq3WrMunMWqVS3nmrUBnzdT4PpBszT/BVA2
3/PaRBYDC8LRsFdrZpzaujJxsnqTDK5HKbJUuoJfGv0yjJubnT+ALNxoPsnxjZAjUrqmeGHFPXF2
GSd5Ja4J+GSRTIR5pvd0G9ssg9BzRBjbqDxExsesNsMAOcv/9QnduuYTCcoKEEZgG3WFgR2X4l66
e8n4GKE1BoB6yxYk/osotv8J2YJWUzU/QsOrRfpnE8eFR8Ai0gS+OCesSU0JKHApoO2sgMaP3cIV
sjbCVK6rQiVNDghKYW3OXk1UtLcg2ro4PhSINI9vWkf7Is9oZ1+kU4t312HDBXVXvo7+kXorXQ7q
dHfjM+O+veNVCJzslRpAOyQbdpLgOGF+NDJMnYT8Y7hKr8A6NpJSCqvYeP702EXfUpSrEYecdzVS
EMx5I9njhpe0GKGONhrvgeEdR0iG/5prEd+EkGfjMU1juxq4xkPiJNklA13PlcLU2forjNX6ZCKY
bNyS1RIZM42STYwi8kBsfy8Szamgj8iDlpzJxzUMKqoWtmYIu8OrTzRuU62ACRszxDE0v/HNyk25
SRR0/dOjus9NQbyXMM9o1XOHAf8RK2tB3F8zkH+mM8oWtEYkNDQ6+6Q7LoLbBkDJXkbFXksxct0v
FZBfvNpx/c+NJWYRIddrDVaZ2okfgqYEAvRFWsLJUJntXUFMJmye5Gf0MzwRYS8N1DeYFmA0zpbO
aaqtjFUOF0pOEGPIBj9TEW8BqhmR+IbcnFbsZE6UF/Lc9x1ZbyfmjiJa40L8NAQQVPNH2jNMjkSE
xiUXigHz5C2UprfXpL41z1UnP3N9PZ611l2Q4la5YTuOhMVy3ManN8Z9+OGZviSIQE24C7cfJIsW
XCPynwz95CvbJUlxPQAP04/w1YLK++/rQpXPmAf5SKj5bWdTpwhRSCnR+ex0Fytu9CN4QRjyYVod
XY4bBbSo38J7MDdZ/VoyyRpS3OjqM9GEyheGfB4l3Yf/lzvCmEvasmUsKXcJvlqL9glyjJoIzkAn
EDGbI8xy8A+5ICxOiF7/B1sKvqcWK3K0SHI2PHsEFpHwPmfrKyqHHV/KnJaeuZS6JaMRR4RKNKTL
wCSt3ylhMjf4q0ep/kqc5pBEDY3pfko1Lf/FQ8nsnnE4yEMajZ6veMmz81fFU8xSr+vrYnzibZ7e
4a91AnbcFDJoJxx7FJHWfeIvLVMbJBUmoKqZGIec8W/Bt0KzkBntNQrf/aXo6bgdAlSVumPj/hIE
VczILxPmql4MLJU9x3z9nGptnRLLOayKQdfgmLtOPm6C52J3o5enz0i1FI2yF1i+AcrswbGbIthv
BxQOZQ8RJ6jMLWN9bWu5zRIzVJK4yaRPp9h+4EpsDPTIcZyK4VQcZdBLBp/2kb1xwbhFdQIr7LR5
evjiEros1DDQb3V1hoROB+U9C0JGGUfxqgKrIBI2ktXp4pR3etMh0e5CTevq7mwXGF1eo9HHtQ/y
+HF7M87RRsCk9je36sx4c2Ko5gUwvfUTtLaoiyHyXUmTZIHzRJvZHGs2GORwWje03LrjwSf2zVKd
p3G+8CTCf2uookcfkHGm7Up72whfX0NdVUCh87KRXu8VXUC0zPgLDKVcU9tPzV8o3KbHx311b1ab
oWzWoEIcmZeA6UN7aQGsZtq/C2Hcq+eD+UhcBS66Q9yPjsDN3waZ49DnYClzXBkEALrGSQy58G2J
HRlms+n5NlBU7gUY+xEc9m3to9v25wSvzcBM4RcASeupBsFFlkOG1bEmVGcVki4Bdw3F1iUx/CQe
bTM5QNIQjZ+er/kEu8nX55moZZfVfr/69W6Pqd0KVGqbESL/coSGrebQqDfFJIBq0RSZDK0NmQz2
57CtOzZkUI9H47cK7O68ferl3jNEpyTJGSAO5fp1HMjnrPp7yCcYbXRomtK4n503tiQhoaGOQgg5
e3l5jQPvgBMTmumOZPzMg6JNVQJhVIVLG+BZIfiNhd/dkPryck9tfFrWjrYfo6/fO2En9qq3+sML
qs++lOlrs1iDivt6hTpNiMqSUInkjveAMH8d4sfXSFO1r+b2PJtJliiP7S6V1nfQyf94iqfcFQPV
hTFRyVUMK0WjxOHNFCGsc7SQ/jmTnNlP8JqythSF31DeXAIiBBWFlBH5pWPaz3nQfwXDyWqizCjL
mdRTlYrYaT86Qw8ayVlbdbVWAhry0FeaqSH6KhQAx7jYTDEE5N9FR5jbNx7icisa0Thaj6aUR3Lt
peP4ZJd0a2T8QtK9m8m+rOcld/VaZhcxrTO3zj9xQuJnVk1kY7y7605sWX0D8KOfbjhakUOuoreo
xfB3lzIieNXwIWtBJdZdDML4HJ/4pU6yOSA+ZkI2j400rpeyDr+oBP0JLrz//5WhlGtQfb1zmWn2
Xjm2RwD7xc/HgEZESqbLpaIF8eb5/AqFu1GPwXKAlBsQgUHBAquOHOfb8cuZ7nHjt1llMaewaWIF
07TYlgi/gWTdezgkqjc8NNhaXDPK43JJfGFwiGYpzHg79B7YfrcYukpPRvGEN1q3C/mf5bl3RfYV
hPzfGOyxDEvgG3VJANJn2HvtSKD+JFqdI27Ax2l1yhAKkBnFpRyl2g6BjOAKl+UrOFTSiZH8Qc7O
+HjZE2RppsP2/b4zc+QjKkeTi8gMSTtR7Du7k3zDwAGW2/L9buDvdchnSSabw7xifRCIMuoGQK5o
IOtEaeYkEs7me+vVR3104ltiFipmio7AelKqZ0s7IWS5qg4fbEJvaZCF1/qC8lrxEXbSitqDYzC5
L3NxvwlohAvJ1schBYaUVVeXHQUdiMMp5W9pfSVvPWKdZxOdbX7bJGDrIZya9EG4x8bReJIW5REN
VXxF1dn7cRQv4hxV7xWchlo4Jm5ES9Hw6H2LcF8RXqUNEOORHSpNNQRKnQeifEDTr0uGGH0zPK5l
sQ+wo8H0WrJgV9Jq4GiG9fcfFHP31R6T9RoRz4zZj/v30QfbsGlsfAfDaLyVPLx7X/BZQvI0NWBn
u3KYxUGgiP8eiRaoCdAC7KOP8UjOJcRNfui9UNrmk4FU0i2UZPUAP7HrnqPfAbagJQnCo5m/JSDU
D3xU3Wsw1J2Srud/5bjXnLd4B7pdquk6YGz9g6ffbvkKPQoJahXdIY88z2U8MuF431UObf/0Luuv
1yXSJcUIvnudMIw+aJnvlPHHI776vyhXdZwC9XsBczevkQqgWIWqpHvtO9vRib2y/j5u9gqWxnbr
ayDp6ho4BXE042Q1DCnGMq+2/nTWw2HSvfphVKMzkHeRuYtNIm2HuTTf/tIRkfxwJhiY5uzkdIGk
xr2Balbw+oQnwjSxE2+ZlWuJQBcvOZ60Hqq7u7EFMGCftnr6CjdluHXdB8Mwep1E25jNS5fZkExQ
JE1Bzn+XGFKyErb4QvZNEN3zMc/0+74u/lAJbQGzj3kitkXA4oKlRkpNRDYwtWuBiaC9YAoC7rVH
FNNy/GorpHYmYIaRvnmlBVrMv7Bsgr8Q3rYJmIzqvkTGcuXPV4lczww1wAZfZMHSjGjBUV60h11X
ozrMgndVLAbcDfhLgFEuU2tLT69yplLN7KQhs2d+BcmZH/mwDQXtxyvXyX3V4MXNbo7hMi8TGOSX
JOF9jwGHKoGfpy5RzdxAqPP8R3tD6LpxpPyJy2EALmdSXstJ7I4mTTVM6bdX5HJ3cHxapugs/zUL
+wE7DT9Kq3qIyhlqU7Uni8mcDVaN7nkJYD0D8NrUpW3Q0+b1iEpY8XaC/hkhffyNFK5cdNUvcin4
rNCITYUZ6gHpTHn0xaESjL/GC3bXCTgEkhbMf3e3tnc9R6PZ201TgZQQ/L/ygAoKmSN88dQmStGa
l7M3eXXp4M5NeoqG/xZBXCWEQudJIL6Y0iIeP/TE4bTPv4U+0lZzgdEmyBabkcNQjbxXWkBaanl/
9nIPllpfBsIO9VGR0jlRpN+gNoSWXuiMgNtk/lXSwmP/Subh9ATqtEDKrD6Ly/FJD9g4rYuHY1WT
NgjAtqGsqlQE0Wzz0hh7ZBYugmeRDPLXXwtWOzWuKkmzP+6nWKj6P+JFfvL/vMffDoowEosC8FjQ
32oZPVlnGFS7y83MrFF/7SKCwvvPRWW8Erfbt759BMOVxDJElXF6vELsgllvQ8enP1CVBX520Dgh
KMssyRIzVxlnnHIU3X2n5qJTA7MWODJMB04Yh6UoauVm7Nqd0HkZQzlur3P8IyNKxKoIYEYSok0g
/GiFWgG4/fnT37Y0KI+7nQRO1fFkhVRh3cOjgKwLzYBnjtu3Z1mu70crq8NeGPDjbhSgI9QKseMa
dGSl5jLuxRPKwlu2R9bXhNSHOpo/lLiz4S3MJNwwyP+bUwsgAhCtmdxLzqGntpwb1UuCElYzoqUC
KCxHqP/fha978VY/mBB/9fI6aTPJSRLLvIFzQ3R+erlvKuOlaTFNpM3au0WacUZ9kAaL/vUa0BtP
lXcXGuNrvW6P8b8PprihAf2IxXWQ4nfvzbq5JnoLbi/1V6UUbtCJ2LoeEQdyGQ18tPUpHtMTmZ/h
RZwhL/ANKvRb0wh+wlOhr6ZfhJGFmzGk1+3w2D9NCl4WLqwusxYgZI9ePsPvB6sLnXQjARZCKASf
5DjZ6EwpOVEH1/oSHsAIOzX7dYPrVQZ4adGI0wlYOKrP6UXBqea+Bewo2Q/Ut30SybkBwBP28d7z
aueRHCfyXJT/oW0nl4AgNTELl/i+fzI221YqKdXhkFHvrfoG4pWrYNUlh5ktYLtCXRaU9SDBpvGP
UowEnvyRDmhJBpt2QCxZAY2K3aHt/zOd/2MsG+BSx48N4Da+YpRkG2nm1RFij4ZA5w72ROoCT7Kk
Z7OWizL85hS8sHzGmKFbLC6qKiqQTd2P2+qtqMGcfNxxAgY5OmgPax7Mmx4c62hbvpzahES34PQa
jCpvUYkAzi0HZZY5uxvSbinfQvqI1Apy5Q2b8ldkWAa8hW6FtYWnJo3PSsRznZXnL1BOJ9KWcu7B
bzqM0HhK4NmbFhTQ1wj88idaYUiDqSA8QtcLKV/S/vXegjWPD/rxyC/9N+EDAfGBbHYpoS0eKYFo
5vXnJ4J+70f7u6hCSlujfU79WLd3WBQubLK1nDfiUOMLVf9x+hatDuF7TCy1vlY4N7Sfq4zahk7b
gildh5jsINbUMhyh5AA6iWJuA7SBqU6qMwZ9/o+lyt9QKOnybpePocv2fTd4sajpgv0uTL4vCkNF
dzpw3Hhmq0vnlVTgx2zzn5h0E8P1VTOuyBUdxUhwEM3R5mNSW/WpoW++/8RZ7/lE1uOo8XkQdOfw
+U3UOHBlO4cRCQZL4VHZzbdyI4VdY6+arZl15jtgxneEgxH14y6mJy1G672z3/Jw2gymmKUA/eQO
5qpuUXXHwW4Xhq19J/5YulB6K7Jr59QbWx5paR5QCsFZFW5eUtTSFDuKuexL1IeGbgwBBh8IZF4U
Efxu1mU50ZMM00TwPi9zSrlHY8W672KOCS3kNSV8EugCJrPBv83Tbwg1bBaEbLZPBN6irSPXyH3u
NG463JVLX1jzGCQH7txPE1lvxSu+lTF+lSSsuM1zb9JPA8Cdam7Mr1kX1oFOplIOEucLYS0dZvKk
3AruXGiLedltra84552eDrLD9FsjzPMicOc7/1SmmMJMvT5mzAQdndnRfJPukD/gAhZXF7ap2u/r
7bB4ipc97Vwb+jpeaRFi6ZzoS+WSz2eyk0b3cnxD3SH7ImlpyTN8fCSc2i9Ft31vIeOlpm+5nsb2
Y4HQEmXTD7SXozUb+P5JqkkLg+GMY/Zr/tKtfd1N8nD7DcBQkowIpl47VrAtRAX0F+E9DccS7faR
X6aCpXv2qmiIeFXJWwxN5gqWiXi62dg2JakhPRXISUj1Mx1DMv6gP8zTv+fb4jXkPIJmMqXZ1+k2
o4BRQYZi7C7uG+KqMgJzzhyHsTdVFNUB+0WUxoPSJ/3SzUdMuLKGEuEROAUqfBvxtfDB2vXBISCd
hx1B1zKF+K/i4xnPIYwOS6VBkl71zyb6jprXZkuCF3LhaPjsCFQwFDu1Wk0FZlWN3mI967R66xfi
z0JtM9fKBWhut2Cu7xKWnhDZQMImI31Hk0ayF85rBg+N/tnwdH+PW1wWxww6QjgZHaUEbz9GzVwm
1oEaaEaPZEP2ihNY7kcLLsLvBx2Qu0AhX8gKAA98MJeBNQ7omIrYqg/yMBIPYxgIV2cnBom9t+QL
WyZJKAzrj2lgXSbQz2pRkOfyqP+hpb66rnjd/YqISRUYWL47YS6eJng6urgjGUbNy+dlMKvojmmr
iMfe74ncEQFWLCxslsh/Yficxrf9qCcmEBikhtrhP4j+s8uSvmRtOykPf6njK/0bLVdxGx2b/vYi
scxn/IALbw/gy77X/MYiUE+V/tpmrp4dx4wiSWNfoGL2XeZ/XSV8eLiBmM5ucgOIs/bWHy7GGrGO
Og0iXqwyWERuOrTHPKRZcJk4im/RV50mlzRwq8Tl0r9Uav0jD6AOU9fEvl337N6OGqAwKVRz1xrW
TTHiefA5ZJyuwQ8GuwUI2leJYLyOLpWLdj/46vAjptih+y0/Qov0A+LufZ+Lez4tZWqHCnDWU4Sf
u6aZJyzSo6QUvCleAFi6KP+ZVuZnd+OOf0DvlFGyMIeirO9DnpObHnfIvKEm35jwE2iurhMZykUb
zknFvnG5jYwBec9FqkFp+2McbDSmL4b6H/tgZ25YTMjZjbJLLUWr65Xt7f4wCyo9/5h30rvo30IU
jaRcYZRn2rME1IV5kDg/uId2rG10DDNLnr2kxV3/EQ+HvJSrOfG6xXJ0xLSNWbyPOQ/njFIsC0mC
0G56DYT5yNJH8nAedYdNpZlHaI+2En/mdwrig7It4m2QfHJAxzLX87/lMgQ2NbhCo9XubUd5MztM
Y9P6DyKCkd26jtQJO77JfkprtO2w8Pdncj9p/CwW2f9o+1UBLRIABxBBR9OFr8dTQsTleyI4WaTl
5/xqKeqC9H/3+BZ0ycymZLh0EJO0mZ/TCaljoyH2DS450PTjH4eXT4pgjEhxL1P0uCXFPY9p9Ov+
YqgtWW9y4XNfdgr79Of0cOdyJWNjM2h0QZfBbkFwlQa9Vw6IGfs+AHf4WaI4lPCADdlxabT2qmLu
2FP2QtWD035pZPni/o2fjNS/XQzdeMMQsLgAmVM5H/OvmV37J3i+lJ/8xUqGTXAszEqEUwaMVL/y
8VFl4APxj/AFOy2N6Q4Fmmdx8qtvIKK14B+Y0fZgsla9kWuTnGcev+fjwiLRmMQrfg+J68QUCn3O
EmEgPkXCJ6rshDb1Tg10IdHPHl7b+LlC9CeE6EsJfEgxtDlnJ4AsGEzCPMNlTDD/GE8iYm050smr
kzjxRMGewD31rSyqsNcd7pAPI8gX45DSQAv3/StgbHF9zMYVh/12hIS5/xdeYGxgpsJrWDGoR4Ud
ki47xTWEJ26eMrGBLzzBm+Ngm/2LE7xOCANZNF2YhyXPfxQpMYiCN7eVLu6b7xOdun2lJNYkJtVD
uKrYDtnd3wxLSEsEUzmSFBoStJG/xsMOmjedRoPcUP37+ll5euilmq42cTcZ8x7PGod+majzPlyR
/4fb6ek0SYQ6hfRPNMK7ZZmeBpzghk67fP9gXJzMmoKNpbsvIuyw9HHcxUbNBxhSFmbquMMwiKPq
mFSa78krQjsb7U1JXMbwq10zEP2iM177YCrxGwqmaldejpgHv0IHHKW18RhFP7E+yK5M4gylmb/6
uVgIVPuvdX70rx4K17+d/AjcBPpJrw3/ys5tePUlctDlQAdbgIiOq/JCOWjDj0t6gIgY+NCBuqCd
XucW3aSGktm5YdDA6wvnclaff9/L6wd7yoAqkthNF9AUP3tsV2xsHdsgn8CAIM+ljW9mI1AooP1m
9I+haRByZg1qhS4BZBInDcyynG9A/g2bum9V2PyJHOXs/kfpMaUtdl+0hVNE/WtHUvWxC4KHsDZj
R4LQ2Z5KQMTIdkyxb5XitJBx4XWABr5qFIDZTvhevIy3yR6unPW/xExtxjhVYS1y9BUj1tnF18lH
jSjtB0mAMD7MDKI9zguIFgIO+72RImdIxu2AyW5gKrMA8OIJk2RCLRC1PU979JM6+2jiaXfrCJ2k
Mc4YnLpR+emkf7v0TKq50Z1iVWFll75zCe/fxVpHOAfbg8DiuYfdtvkrURnVSSnHNoBqxHxdrEJ7
iCMCoMe44AnrYE+42lVZR32B1CdD04OKFP4eDzinWgtG3N4grtkOY9YEUG16vYwnOAgulV/47w5B
/+k7kKh5kBm7f3RF9KPoMRh5uxUtr39sIE5DEf+LGgbu03MXSpHppDqzpIsgaSmbhLYuEBqc7okm
uQFbAncWE00bEA39yzm5M7uwywmeMyrwNye9pb8J9AGK7U/gk3WTAzqEBfvy9zX7Xdsn97aHf8T5
jJbmLtJ72Uxo/Ri+SuA3Ublki4ETB2hnw7JuHQVc1gNLES6EZ8oaEFdIJ11+YJY0Hf/FrACFdLn8
D3kr9Z53o0VoKHO/3TYtWvO6mP4Xm8l2VuW/3eXFdh0bLGA2RnawxPS+2qaDxCEe8GKBJAzAti4U
Whhbpiyk/pjoYiFe4A8O2MT4+yHJR6U30K/NAqc2sRBSmZxBbl26wty1Ya8HsCxiwCBbu2Y+Uo3C
7raid599yGLp0AI4oXJIR8V49VInU3YduAVj6PuzeGkG5Bh4i4OKnw6wosPjLX4et0MSBDSrB+/F
hySra9ubiFx/O/XbSuPApgRgmRWnbww40omUq8axU0hdWTMwsujCNZ9qbl6U9iExjkgp7OgqApSd
IY2TNhalCmO4MGDpmQo/3LwW2tSEQiMthoMj5gEJ6cMtuj2L18yzNbKaGl0CQs9xynV7RArGYtZv
y6LNQHwcDO5cMcWAZXUA+0zUWkjDI4euY8g4RyALJ7jL5OnNtQeFyP/rnWrlHCkNYt64CxubHUdz
Q9/Bj4l5xKAB2yuVOZSwc3A34cu7H8wbmzhJzIu8AiVwXwJunF8KyHY0VpM9h4wp2B56dFC/krMP
N00z/XLY/uk2/u6Hdmi5/3UBREoRL+E6U1ZI0RX0TWwPPTVeP/fwVEBavZSfkisktqKSdj/vuAqh
kFkCITAupRKaeyOSTk6zS2HLYJsn0rIh23zXotlJdXrE/Ls/4unvmC9/l6475cRMJmfgis/LR5KE
c+Via+cw8/lZfabjsiqndE3DPhlusFw8ZTgm4RGxIlF7jOZS9QbLQ/aUk/UElaEGOtDZR4i9hN+M
aNaZ7hMKQJdV+xYyDNT+neJcVDpS8WddX8ZsBJsG1NApcZCzMUtcagBq658Z0CVaHoK9vhta3j/9
ahDcvEpGq6WpXdGWYNeq8yHjVUHzNu45K3TUDLp0gtdvUi1eGuCdj45SEU30fyd/H3eMfHnglKQi
jnSYCPnG1wrfM+T7JSv1hxs1/vmdzJjuPbhhLLelv9kGu6Opl85/pstWqO+EtBgcA6az+RtB5cUG
FIS2IdBbEiNFm6eVrASMIodrHCvl23Hy0TJEZ6bYMJT63HRGTAIeYvRoC4YWW1Vw0aYOlk4dLPSm
cj3irrV4TuZrFbvXCH3EGmTW15/AHBBHBvq+yk3LyBJeXYjOhQx4RcZrO05atIW3xEZTqDWgBcmD
Av9AM9gOlNIw71M/eSe1OzFd51N09Y5yRcCrWZANM3pA4T5/7zIrKLMfDMWkOWCMWxHRtBwPTLZG
Dummt8VtL6wkUbgBSpK6keQ9Kp8781uJHJw5OSxxk5Chunjt/i0VTQ/YHsYPAaxRd4ck86Hg1kWm
NYiOqLojpyi/IGFXoOY0b0yFpoE9NCeJXKBNFYv0NYc0dvhu0mZc2lphe08/OIp30TKrP/mTOWx6
WfYnyNNTfgx7RHTW0+VuOZ8qWuKBBX83s0cUI1nntxIiwYObNyw2hqckTUkU75ge48D5uNNP4JS/
NtskKBFGeJ1CV8Dseo7sC6SVhWrJ21AutJIDgH5YuPycCZTkHgUfLCwD3m0Iu2tRdt97O49/3uj1
1XRMoPKDB0t6xq5ODIkxGZPyEBNGYZ3bND90M+oZPVeiZSxXIpbc3eOhuv3DWoFKLy2XYv8AGjaH
DuGZ3NiZc9Arbfnc0pIkgdeiTP5OtPO5iEQbrOMvNbhOLuwMZcSWJnEjTp72Mqqb4R2ULCWlPTd0
rEY2vMvvv7pO2ww2m4Meg/3DDRM/NmO0VB36q4irDE7aqjQNJeXPsyffSpvQablevpVbh0vlJZhp
/qZDLPRTWrBnI6R0O5DFeTfLjmZ/nnDA8v897kW9jAr6SMlNC/w34FaCzVdDz0KRycmpDJkWtHe/
jgioYCujECVR3PuD/kDVzUMbuvIaV2uoag4Wm6sArK5Tgm5kBJWG1pSRIPPFHre1b2YeMXc6gj4I
F6ZLS5U81fDgcyNvXoANazVE/QikhhWpnzOlWz+Zm5R73DCHl0EzTj/dkgZ5ZEkaYi2lxdm/5sP3
sYu0/VJUMPitzv67/fAB3G5PQxVFy83OYeccKBVL2eoOQ6cfYYR9w0K5h9fq9Ccd9YhiBq4pnxFM
QzosFTHd6SZemMfkRDfc85JINsyarl2iIsQ9r1MzYRWXcjdx/vZ8YLkQTzczQgJXRkg2mjlHttPs
KnuUu2c8Iv4r0tCX5JLd48S5No2RPix1RP/79lAkhbCgY6YgjmGP9yZWfX8YmPIT3+J3vzJKqMaz
+RNAoJW2ohyqsoMd6R+xwzKjvca5162uJtLl9RQ43tUoXZF1o4wmI9nvg+b7LhPbf3onWu1L2vxv
ffYzuh3wLFGzuN8PRazJxdOXLIslvp2cn6tCsKvj8TjlDZ02UJMJjaUwDDGVz6NLXytUSQEn1iDo
PmVp5e5snJ+wSg8nyiFXJvtT/J28xM+SDAujWN54VGqzPi3h7NQmgiv6EfxBRv0sb5xNLyKvYRza
SkapxB6YQu4cMyU2kG7b3bRfNRDx2JXCh9ZDnj9XPNKdu2ecK3HdcmecEo+ww8b/jwsohgxAWDXz
GBOi6HZgqCBNjuFq+Ykl6DWm7OtpbD29M2QJGPXbASoLQsf4SQKF1hGpAQ2plcumqzbkVTCRy5mF
X+HqbOULzdysE12VKmvIHKZK00zqVxm98V7XC0kYwFRGJy6qhEHUNxlCzEPujJcO7tCWXEOvOuL6
nMYNjKVwrx8iq1rhaiUzqfKGgyYCTEVHRpERxl4D1ETPCrG6lgHObXuN3rAJMYl8RPJLRQl/XNgI
HcWWBZ/sj+AMvTJuBYxEmeVtx/rKCTtlCCKTKmouKIeROQD/5n7Hu2E1f5Zr7zcjgPYcyq5aeaTE
hrS55+E2YstqJrI8Y/B9Dxog/i9mM7u7JZmJsXGukU1xla/jQvUH9y/rLG95Cw35loFWyP09i887
a90DVBg8u5tcLPg6+JtRG2oYvmfUgg3LyWXqDALoXvtX4FSVSU322RxUbIcvB2VjCKr3saJNo24T
7wdvRGejYrymOeVgp36feM3De5ropU/XW601ZM+/vkZPJ+MBHPZv/BeKrYWkqUS/h8gbmcjk3wg6
Ekb+UJxNdFtqUBBLAT7PgUyHEAwgwdMFs71pORZP/35zpP2/HkZW6vUp2PhTR9upMD0gEadT4D4k
r5Q0w/WKgF223iyi+4oKntGtwK6OK0jswxrwjgVrr9o0TpjhQnWz5CsD0bCLIALO5UIodhFDTO92
wnhQkbH37EFM8OA0HUSMo22ViZqtVTO/BUPNVx0Z5Cg+KvGPcR3pPSOQ+ddo3g5l5KWRRBkKhBQ8
Aw6Itl6I4IPhtNg364sAZDTI01fjqgeQ1RR9ncOEkyM93n5WPkZ6gojTOzeEO5ta4Qe4/+QFscNv
mEBLvWzSjTERjVD92xgoI+ekFRA5m/j2Rkv9y/T9XKEDLVRChhPzJa+fqcPNOabxCefPAGt26jKt
LqeMQHoFwNzRcncUx5L7Ys3/OiqTxTcar0AhpFJrbwHLtbs2BQYzrcqU540kIVRVlCH6O/jYhxwh
jAvzL8wur3Q1WnNtdRX+VdQTb8z3AWjmX0XVze8/YvL1GlkaZ+5mSQu/cgPO3WeRYbyW3zFw++zM
oQE8MoLhA0vpGaPVmWDMoVGTBO8GE9F0I8UplDwlDrI7qYG8n5kKwprYgDITUYrnlAAtE4m1BjaT
U60eTzSwA/kNx8yTc6X7PEGSuR3FECiMLryTQK8nVgVATLIO5eF3DeYGzP3NrzkRxXIxbpkkKibO
5/PDczdMkGcZD62d+O+wXhM0zS0ZiJKa6FJTZ66mh6+EWNPx/M5BXfa6KTaDY7H/1RnIluTHNVlP
M8Rgg57pYwitmH4OeExVdQYoAuvoH200753cw5Fb0Wlq7BJUF5+YvUh7txN1h0ynhHT6Digx9uo/
+AbyzpXVqN2+clVjZXlEUEpDRTRj0aUWOR4vsfl0/k5KV/LAPrdUwJs8pszdElzSExPRSSudU1Tx
pc4G2HUEc8xrNHrEtR4LtjkPRkI96sY8x1zyBCt4w9YIeFKNWJzSm7JlqbG+U0xNZShBfklb9rTJ
8VOPrdj31Q0lBzuWI8eu4jiuLFqPUxNooyCq1tJF1EVxWBTypImKwdmsBqxPWLPtiaWA6GOk5t5x
69vYC0D1X2DppJocwIjRN9Uaar7U6WJLvd63frCGuNrVnFl8SuCqjfk1MQZKJYekrJ0khjDFoSGh
2FnR2mGwKmQPtMxPAbAHusi98YjKWKKGD9LOZVyln+2Vz2FKgRZbKOSQM8EW21bAD/C0LkF2hpfr
WJWv8c+0mz1M5RbsDV6eJzRaERG4yNvBOBJoIiwMOfyZPyaSy4eHfrxSunfbijdvnv/RvEhYNRev
RuCC9Gh/PxN4U/yEgA/55Sv6zCz1jLJOVtAn92Fp4jDKsXMOckBDHWJdXGhCcOmiokV9fBQVud7B
uOJ7KCNd1TlOXcb7NHmKUh3fkGC4z9pXJU0AptUwlJu+I0ipKsavXibQjKGWmTGIpdQl1KSmtxNc
7K8FRcTm4V6dGAZg+Nb+xCpZdINOtUBgiG7IKhh1BGsedK1r35qtJbXiRhYDJlzAmnlOvPmrKbgY
w2uVH6zbvYowb8TIz6f43KQezZivcIrYu5t0iNLizV9cwUT3arjGjBuX2GpJxWOVz6iCMm7Vxceu
ZTsg6mSr2r7asbe0lPC5wiGRSUjrcB9K9hUMVckgXux/Ul4iE11BsqdBGmzk3++37x78NI63LYHB
ZBF8DktWn8DBLiN0OQAefz6kbyr02U9Xc3WyrFOLi+3b2F4lasos1ui2iT97Da1vnxbKZGs9csdP
THV/b/M0kJQb3ImkFCIzHbfbZIMxTutgjhjhpKcU/NyaWrRfbORjIAj8dob4bbLNS+eFr4GkSLRi
/GG5kdu0zJPpLkgXMTMm+wj7XEey8dgbygjiSf7GdMnKix/BGYgmHKy2WXRdTvhga5j+eZNWdHrV
et3uSXY5iQ+cDMEZH0+892kWuAEVl0x04ZziRwxW0bQgfU69HD7huS29ynJTxorcFc39eaypuQhz
F4DS5nO+VIA78h/d5JqI55OV3WyxSeL7DD4xWP0DULT+I/hErpPbSwlyd2MNsvKAtH5VU+C7k2x3
izak5jofMBR4OjaWwjrhYaIRK1OsFtFMCETXDImOigu3jQmC9be7QjPB+lBrxcDI4VaX3AhqS7sl
SmDUrl7s23RqZ8vHo3/3AZ5rCAlVUVi2mAdOhaVECRJiNFy0TFJugS2UkA1bYeXC1sbB21x2BVkM
0h8Q7iIbwO6NbkFRt/79/gernaSnKFcF6gTgnA4EhNgXcu2I3PpH/1LUI/QkvQZH9aIOUx+rrGus
Egde66CsIgxgdRZ4hu9gpB6VGgFAb6GDcOIux1g9ARg5rkk6edDQW66PcRQ8oEUugebxk4tZwnP3
lyMv4Z3b+ZsZbKTqjjnIyHIReMzBJHmmvM2ZdmlxaagPR60s76Dop3x2w36BhxMavoYw0fbybtHI
gvrO2nBAHUmbYHVF3/+T+PRNvMVz6Gf0xsbuXcxzzc4P7x2+LYGYI3Gw3AjkUm3NJKoNg3rqukNJ
UlFgZCuzrYbi93rPiYa2TCyZrYKUung+D6f+XLvDnjRbCNrg3MKnfDKPXv1dNMeGVL8Wc1e43wZV
5GpPwJfU/XbXK2YF/W1wLG86iS7dqqL21JF8TQs2/gts1dESgsWRl+mgbOxZszbgEC7zs/m3wqsn
zPbpbu2ZLlIxCU6DI/tpDx30Kv97AQ8SAQRMdG+MBNs3M8PO9nppt1k/4E1TghrObX6RxQ23SP4N
rYqsRSLB5M3bTPmVDKgPoX3qJiX9JSbSz94hFlN19kJ4NXDkkIdbUX45uDll8B2qLea/KSw4AeFu
IKkgITMj0NtCVfzpdOQwLRDnp8k+1SGX9DAxaspzCmh84qko/i8mYAE4UsK7Eyv83UwNg6MkZ9TN
r3aFLWeQJuDo32ZIcqDTpBCrbLUPAd/hpv5KxmDmDyW1Sv2MKEHrO1334PmNrBc3Jpt5C4k8aPpp
UkL0GkZl8A1xpAWxWzjZbjSbkVR8BYHWBGE0kr0cFYq06i/YWp2/wo4NnfPeWk15tw2cYonQ7QKt
pzVMF6SkpcY2RdxZaOgndU1tvM6D6u7cYoQ6QzgCLNgfz6k26OAaqit7b8mk95+3cFo2nIBqRTj1
jyo44BPBWYKFUbTXrgo9w99GWnfD7MTV2O/1UVHBzNQqtLjnCFqIsruGd6xDEV75h5XPOdCPK6Mg
/Ezr3eo7klKZsEkSPS65McpxcPOjitGCWtoTuCN2OdRlcQaTpVBbBWbBilCYyR06wyuUQHneIoUa
5rzoajNECfIW8xQZk4+OFabM42MPmifJBmhFWhrdpdzcTsR5maA7Q8h5/gfcNgoabg4MTkIRBC/e
lYJGpu5DWz0ex1KZ+cKK7qJXb/VDeIhfwtIz6Eh/9mEMnGhtgc4Zr3M5jrn8YDKKIOi3BCun9Be1
/DGBlf9p6jLVHqCT68ALEohjnlM99mVuqs+h3PDzMua8if/e6uiCAF7/jcdMwrJF488lbc1SGhvQ
vfvF6+KDNH63TCK7mT5iPim25AxCDfQIdyKQgkSEq98v8bnXMMUoUwiM3/B1uOrrRaRScFRYeuym
VTFAMbbB3zLPT1T4ayAV0oyxfR+4c3qIrHsAOalonyiZdgEoojHmIKxKlnwmTgvS7BTzqlB9pZvO
yFrin/PsEark0fu5qA9y8mwttrtQPE6MuWl4ziljOi3T24ut8er7Oq/x84ydjQvmiv13RHya/pfq
ITgG66WH1UgH3Gzl76dpZoIPrmIkN4IWOiPgSWzh09i7xyNNGFL9S8WdzeirY2w/DdNCFohblUbw
y2WgrW3Jw+vDcZ8JyAFMZZ76uWyzoly8yVfWuH3RblReZk3zJoWHRLuAvufLBdvBGgjCBRFg1q9p
uxebyJ/o6dLizdkGHbjtM9IpBhuHqFK7155CiEycJFnrnELhSzACOy9TsUtqSfNeB8AikifB5cgJ
4b3ET5a7Pwv1HDRwZvPG39lbopx9QlZ+c2BkpFJzHzj9MT5RqQDXY3mIRHNMhfwBeD+czAX1qqU4
wSWgbWn0WRTECuUHTpjU/RC7CJfq8Y9n9aVghsISFhXGd9LOR9SVaZQJUI+QZUPenzRG/lhsAIY8
7xlIoPWXmWPIqAgU2Q6sDG/z4jZwhG+qbo/bdXjD+aq2FXPlyUNvuFWNi1NWO8FVrDQeNEQsfCIX
hM3KmLcbK9WpdFzCS6ur4eW/oSYZLnvZAl36CR84vAX/SyfZfxuidHc96D2smREJ8mcQ1ABPcF62
/J1m7v43XABDylBOU6SIH7vGuxIH2IJz/F6H2fWwgW1ZsCKQkF9pRl9O8GoFxQmO0ouqZyHvOU+Y
QxHUnzVIVx01Aq1S85x6eMMBLwqIQwiidnr/wbHPFHPjwSaSyCIvLHlscvSiR83O6tld82D3mkhV
cjSaBP6GQWKgYt+oEye1QW51rQe2zURUAlMFA139KN2MoghuuXOnV65AUX343Flb8ZQsF76iLdPW
e4GqgBAa1Q5SGUDgxtac59YDuLxen38K9pSoM9OsDGbqz/G2oVjkr1nZW3R3eGTtxbL1spF97lYY
93MM7gnMxfNT1MUgl/ESdKU1GMmO0f3LypSYRkVmpeaKQSJt1s0KX3fU8mwFM64zt/xiwIWSwZi1
74++yAF+9tmtlYcMsAHRt0tpeVj+QIJBnx20OIi5A43XjLDPqqZVXbgodR/ntVRxnVcVzj9sz42I
WO+pz2L0TtMWTGOOaSt/IErlMLKC8vGbnttoWU5fEVIxosPdWYxOUT4SrmHIW06K87Nr5g+IhtrS
K/E4hylzSmR4+tw+TxzFcorDVbz6ASCr8KnaPW3pSVx5DVEdGEwZ/kDt8C5jwCGq1Tv+qMJLdGEc
f71uS3p0PKVEYaJEZwwoH/KmhQFZvc4FIhassGz/+4A30vUZXRYU1M+DTWnwJhfcs9Ycc7bm9u6e
6hXN1zpsBtlxVPjhvbPy4BR9a5boKRLPv3HcFQjaOUbF8NzRX/E3dtT45StCc1USD76c/vge1iL8
rFAwYaLwMoPVY4Ftg/uBDFjwthdTIUaPjF0djtMWcVxa4C3P19jlqK7WFjSNjQshVUvGMIKIW4Gr
QesJcEQ9Zc1GbCCPLcWZiJW1GE4mmvDPtcscrekq9Lg59Pl1Rzm6/ROwsyzyNzoecFWJTKO4ZIbT
sJQ/eSu4tXC9TPgdWt/2G937/wE3zrgMiY3n0nvEzS2eSu+3McMREm0jeXBfUgChn0MrKgSwN7xw
q1ASfC80BOHruhfDWCPjUNm0qJz2QV2Ui5Om2XEUf44ZPBVEcaO8+Yjb/ppyYzXu9T45Mkwa0tcp
CA2ivtBxowBOKw1r6KNzxqozR2S9Zi96+oHB/mhTwoip1ZjMjenWUC9G5Wl3nVNc6fPNxzXrc0rO
Umevk7dipVWJH9IlGEN63yf9aAf98kwcWePC9W35T3CPWyQKLNJV2Psr7Xj3sytJdtkHNEkkZvwb
ayU2AEDacEOjMlIOT5h4ekYWKEY0PuxG8HEsSyTNaGPMc0bzU95weikmwUTWpzheAeMqa0X4MtTp
nD3TwRPZyAVmReY8atiZjkchmM0w1Ipq0SMpJdg0uGDJ4frJgcis0Bpvq5c99BRZQxV2n9bXfReA
R4xjTyJv9zdcganZb0gYncxMW3mqx7cpwgqWYF/oO4c21a4ts6OsOO2kWZznRUP2hXWLMPj02tJV
z9chw8QGXMAPcE6Y8jT5/RtfNNoM9xME3D/c9hQO3xcAuKZ/f26H6DjtnJRRIo7b8RZi4z6U9AX6
LABz/I7n0Igc9YoS9ydiYDO20PHhcfMJCJ9HyycCSCqymS2+nCWl+NkQq8eajhPXbQPy019bx1Xq
ZvNbnqQO9NrCebaX4UDgGgIh1/zLJTNGCFvDVcwNKC9+qA9H+G8SKUmrjVGV2oXRqR8a7D24+4xS
FRmIO1v+hJBCXRPYlBNcN+ijNoNgBl9Xw1OwnTE7PEJNf38veWDRQuHPhrmxOjWsu7T9gc+xAjK9
buA50E3vqVzQbhE3trDhg4tvs7+onvhGmkSIMVd5Oq9Jw9w10J16LTrVDGuQn0bGC9wdK5Ob5ZUT
EtSwNNyY9mZeJC87xb/1PAidkmkEaGMl+v++LbcSKcVw20BfhnGpjhtOMolHhqXGjXg+JwaDlw4J
dsZbGrRZ/cOPbGgpKfOjfzpHJ8cKRghYG0lOuZwxkid1hKD0zDDVxWP0VUThSRL2HgOV61+vzSTD
ZgIKcxM7aYlNg0fQbKsnFNOeHlTXoGsot6YA2Nv7pdzZwp3v4fuA5uvrkhkPxHC2F/gdg0Q81eHO
9hH/v6k8HrtPPHLOBm3IDLO9LXXSAh/lS+EafNWAA/VyPA+26sl51ZxJZ89ONsFcEoQO4y6i9gWh
RiusD3lAk4g3EbqqBX8dPSAUlp+lAO+pyvjMq4mBFdsCGwS+ovNeRP4T5xW4CTysFS5SfMdmKXvL
EqyCMJkitTRj0ngYGMdst046Y4WmTc5tXUBAt1zgdHMJwsCgwpGN547AJXRLMs32o1AEGPcCZuVb
2M5tBwsoMgtIjMPiOZcX4ggyGu6UxA5wGvnpy5lB/dc2R/G040PC512bxWJDFZM0/w8KW0ljjBKX
jvbZj1nvNqQOgUtOvfPXEPwJs5DpkJzUQvT3hYlUoH47XCuX8WK83gyt5fv26e2QxZSPATWge15R
8eDNMurgVIh/4iNf/dqd3c2gTPwf5N+o25NOVYGc+9nJDDZmcH0G2JlTDl9qUeD/9UH1x2jNAAAY
3h6kkBof7wGcoonM4xgd+G3Mhgf53jGfFHmuiu4Jj/eVUqmfO/AqaLZgvihZf++G66tLTLKcfljo
/wC1ePO2A2qbo9GQEBezxE6PkwFt4nF6rrlinTNOH7wwfhdSX3QR/EMzh6BEMI/V84wz0AbK2SRC
IcuEFTsHOhVxPTqZ9otOy4OTUzzob8vVS0iW5ixQ6NmDiTMHeuMqErkN8a966tf2RKyshJaCh35Z
LyehFDDJPJQ941FkI0zM25HX/L5JfjeXjFpxwIjSS1wiXloS5Q7Jz0GwhXoI6kcBZ+hpuOToOL2F
HIQ1Q34UirMeJ0I3SfXW6qD8Tx1fr9V6aaQqCNwGTudCtdjAORYxGDt4YLsO4FSbGuVxKbUBSZ7X
LvjL1xJVYR2+BXrEmd34VqEvMXA+D+mPvyvXCMqYvS3U38D0tKrIHu4Ehjp+6FqnSmr4PQ+P/Kb6
TPP8BiovadCbBeramJN3ggYG56+Ck5KNk0TzlLNE/hCZ1rcLSOP06aYMT1qOWOt7zIr/g1B6ykId
DW/KE9n7xKh0lg2OXGZesTgp2pil2IQTur9jsN9DkuHUIO05S8Z7ymx4lIzVeD+iQ76a/dOMOH2o
OcHwYDpy+ysbiTg8Vy/Erll6AEijprWcfWkvSS1JhQpVq4zLcmG1VBtmvRz6hyRIdMhHTKVZKua0
C4Udcmmt0Eu5LSxPL03xqTAuiNQffnNfzCk2n+RSuUC8OB5rZa+FXI7MI2hq+WrAwHLTAiwozbJ4
Zhr+MV0qEv9xJq7zX9Mr2bFnAwLkiQ0O2IrasiaseqM/kQdJpCM1RCXF02WHyZZ3FD3ZVXcOQXZV
L4FVdOTPUovK5vWvKs6/2TyJ6FFXhhoCc9t4IW20x10fVz1s1h0E4xGmO0pG1DchDgpJkCqJjHCR
TJz/k8sg5Qi5dCJE2vtJirknEq4r04rIsbvGkm1HWuuz8KWGegWYAOdgpevwHr8Oeyl3axa1OhHg
cN5kFXBww4IH6Ff4Podd9EIg9WiwwZYfIhYSOOQjGzglvt038kKNdwzI/Fa41MD9wR7By+qNcuyd
iKsWvibUFM7ZOYUyZvOinEi3daAmDqLSHYqASYL9PxvlARxRdfixuEAr427LKwV6+RAsMVS+fexU
FejBcdM0ERWVX6pIPE3nVnIg1pRTLhA7jVqMwmnaVpgMyO94h5Q3nNkaTU4Yn0pF9R+oeorwBwR9
Fnnk6ohG7rZmT3JCbeZiGYit5+OcT/NveCXEVGzFlQQQVwLl4WGT90qKaLT5ZFDthiTynXkxssFY
ts+5lvyL5h7OT5zkAYpPcysm/YvLSelAfJ1uic+k9XuHN94y1gQWo4/DgsZvHuqaCWaDjQNWt4uw
JsoRCHjeWnmjRlqfFUskASCfCObYU8QWGzBWfnW8xqhjDr13qDUycPw6r2dYoKJb3tkJ9T1xndid
2ZVHL/h6oXFpL/DMwySE1048nY3Mc97DlL5CMAzrab1Ic8u8oAASwoTlwu9N1CRQ8RlztUnfKIdu
7oTpcGdoUnaDE01NS1A6EdLevXVXXWGkMiB42wrvBQsyEfW6VkMO7NknneL34JzJfRLYOCtswxoK
PYmKtnO0UR5aCelsY3SoO2J4+IWDFcuAYm8o/zPNTnRfIvVUe9iK/RDKynP9PIrfpttqW7zochBa
nRaS+qcWY88+cl6QldCa9ho+71TNctJbqncouRQ80kjH/QRjmXM2QfhHtCLxMxj4nD9vigGLoGko
KVcDhhr8xPK1DfMu2CKaiwk7+mxoifq9OsYbu79dgLfHpk4XjSc7Man95wUfvwlgX5/yAY3QUzew
g7dbXbPZkx3JBjieCM4HlQAnD+TTPO/9NmWRZi/IifuAr/GQDliyEdsZOleJIMjYTh2RSFAggUxc
U4PgCDdgWr0aRgoRiJbksT4Nid67is9Ua/4l2MNUzMOVS/zSH5Sd7tT1/ypqtcxgPOjRFqIyQ9ud
1lDWx/3D1pIKdWbTImkfJNGiK1NPP1ZyO/Rkv2otPyjcY08F38EL1DK0pzp/05E7w8+05XaBxLVs
K7qhi8POscuSiMqe1weMRPYinjR/7fArwSAk3KK5SQs6UZDO2zOykWn/9Dv3JhRS+ERSwk00RdVp
dKcJBGnwNIttf7m8+Ll/sF1PU8y56Xv0ZNz0Sw+gzMFbHKdVcPK1WjR7sG0uLziZOqkVLTgnhtIb
Qwju/5SVZJ6KNCIfWniJOdBmFHTrWHFhN68DHdun7adBrq8iPZDHeFjyNb33FIC+FMeVmvml05D6
JJGX/rSnoxGj7dJz8eYtgu2GaLFWkVbMHOfXLmWww8KTZX36fGghUDl5I2QF7Sl1aI5S3KAauOzW
MHerg8QP7HtaS2PJF4eFHOz9wwMmOm41kWzzfhUwiC8asVn6k/mFh6Za6DoEfPtP0+x04KecA0mE
C1t4hqicWb7MRB8O4M7DeehYoCnviaxe6GeKSf4z7pgY7RnDJD0GJcIOCuHLWkqYwRsunltP5hxQ
nM9XvtaDQMhCx1jttlJWz/8gAe3GvN4KCmifIuvBK4Jem9N6q38lqQ+lbwgc2iccpfePJo+QzK7T
dGkey5QuzbVEz0gyA2/+Fe99opSFFDWdEpwYFEVuP2r9G9zzlLBlDa18aHLff0Ix65rw1zmQ7/KE
teRSX4P6Z9dLWZjpwxfC70UJ6L+g+fbnacgGoKzSlmT7ME2rpa287N8anGhy7mxo1K2wjSBHGGId
1oFDptoHW+M6tEDl1TBZkjeWhqxoN7kM35wPs5oUie/W6vHqkZbcaC+RKMVcfhPBNimoCbZ/DPsP
HFrFqphfBOKWw2LlAjs3eOc0YXtuDTSqDqNHltQ9KKg+tJIvBBTJBCtSA+QgPvwSbTCYXEBvaxPq
nfwFA08tOmgCHLWSqDuZ7xypypkRmBzIz7FHopypaex3gywdA+Sotbw5AymnnJXYMfb1SD0je+G+
yYpXcGRKNupynAlbdXcIVkvtIPfbY0tg/CV8g3udCporUVbP7u9PJRzlDBtv3N9Ce0E1qtZfULs3
knf2TxygWb7WdG/xXiTPzqMu3q4/TSYPldbpevVD10ws/+oKXV9fnvU9sO2TeKct81Ukat4f/J5P
9b8755pK6SIZqNO2/BBK/JIc4t/nxk91VjUYanjY3ItjgqHUaMd/u9VX2EETpbA1pVivNXIFehXJ
GlOg2322zo6hW9TKYNmOPkh4IZObqNPDEh3GRO4NDKYMLvtf/WTAp4Ane6hTr5qqwmUlw9xCVdXG
AGWQTcgwbIJlH2CTDvpOOXAnGBe8BSCTMK8iIjBzvJUUMP0nniQxfVZjxTrJTui5vtbxSC62C7ie
sYBionqgfmdGVtOYEscYqiRtTaPw+nml21gKD9GI2PyYSdYD5Tn1SolhTtbohK8rSOWoIaOsxBVu
c+Qn3C38gb09qF2C03kv+MV4YEcpOn16S1iC1um2zpjnBtXNB2va+/FPzcp07qxFlsX+Ksve+rS0
baECKoHVCVVCi4BFV6EAsIRp3gfOWgzJInuCfd4XMI0NRJap4yOcqpi5fTVN97ph5EEOo4XmOeq0
pW3MMXdfPFugS86j/wGG1oMng5RLp3VUTRngTZLlqsB7j+65UOMxa4QthGRWHNdqolHqWJzo7nUP
SMpbXxmGlvndDXvzFxA2eXzcyo7nhhAxK4p64jsbK6NrDGNDezXh4sXHeGZcZY7XeCQj+T5ucxX3
pr0nTHYh2/cajoPhlPyoQQVFwYpKkvgCqIozsGpQSseZxr2hC0Hfz8WaNwGf14w8/FcntV8hRJCc
5JY4BJxMGpCHPzw4zz6otwf+co/uFUobXT7yzaWk2e2mFEuG9ZOjuDEtkOKopfo43vrcmgBCMvFX
1F/avZjuxuTvZiDcfOyOBLbadCgI2t+ox8q3+fYFTblUwkfzoQkemUDgvzqqq1j5P1lgsx45lZ5R
GShK8h3bsydo9KAdrff6VapRnl1V4B6OluFgV/ZYUF4ZLatnqcKWanPURCBQrHVtQtsDDmhyFVU6
pJamm3H3JmFTVYMWL4O7wZC58ZLdN6ypTPvwfaAFXfBcavOOIMMnXD1k8tStwlsOG1ZwZ4TAzLbE
rxc4NSZ7e9TVHX6jHbu66c8sbkRdHBE44Y0YwEcwG+jq1JQhj6SZuXrTKkfZkwB7SZyqO0Gn6uaH
i4rS+Wz+njpGX2lHmc/P/fktkC4V3ujLzq6BfwOoAOh8wa9XsKo/391kY6Cmbp3eNbTitrDzQlIa
i89S4n5ny3oQxidTqnpLyPEj73lfqMVnDTMo7cOh+rHnk9oFful8Yv1cGxrEBMeQ0dApdu9FEHN9
0HoRIf469vobHrDHoqSt6M0m957XlMZbjArkGpRzs03mD4RAt6Me67/5cV55jDHMJfY7tQhgAZYQ
JlnSpWrnB7AHQxrSzQMCH8GcOwAn4k6shaIlAV6yOI5DyJYo8K4g882y8zAVNeqwKNEwsp/AbyxI
eUW4DAy5VdNYppFzMvI0wIMYEW+2m8X1WG5hSdrjT9sBBD8smgRSrPLheh6l/uAkXupNg2LOXeIZ
erVeJuCLA38mMTFJM9glX06O+SUBSShRGCf7dZBQnPPnMdvN0SEeNJzgIq9Loib2jtwJ951QsiK8
ZI/m7vI14iE3Pslz2V1ujKjpsOKQ+ae7WIp6nXfk5vyY4rXHHbGrkOI1ixwHR2PeSiVFhCHuS1Qv
2j224TP+nT28REIKmr5CD3/GHMXL3OF7xe2qgz+wS2c6MYmJP58+XoptHY5JJM6VcnsJQQPFkw6u
p1JCm/KiCAsk5eszML+Ym5lysxzYymMFiDQT76sA2haAybUbr7W+qG7yw6a4k0MeOD2PRWIRStII
bfC+RPcM053wtR7QByT6gzTbhhSvRmSOfMY2sz3F5cMmT0lZ2myjoArxaCF0b1vKIEk7xYy48a16
Ge8E5phXMRGI8MYO2N/SfMSdGOx1c8Bo3/fFqZwJfFZ5XlXMmbCow7DYK1q+P9qJzrwR/dJGEE1n
uQFKJ9NPRnN4yh496rcN5LWgFiV5K9UNZ/V5rGwRWa4mGrt2jlQJpuYBUV2xCM3qQjxeMtLSbJZa
j67ZuQEB3JSTFho3Ars+59eWUoXpypI7DPjJ+IufqkPUo2LhPsNXWEjgIhWhq7tlFP/45gXdaxsF
g4mUK/C0VBpiw31GBV3qqwxzUNAWVW9BhpD5APCWfudEoxvUZv7A8mY2MEHZbceRKtZICV0+3vep
j1+R2hpBf+wSz3txDPdHC2yWMrNM8xSc39mHdWxtgSk43lxc+UEmLkoGCopC2896ewrkkyVgfIv5
hYJo/40tEpy1bYgZwT47ReOTWsXDdAUUVpzTrnfSfD+Km41nKlr6XK0QQiet5V2EI8P4k7Bt1tKn
znaoNgSe5Uamkr7rw2nxSBH4cqLYpn6Uei8/VsXhg/GZtXcKhNVrlwF3SBFLVhR+IelaeFGnUku3
H7KwWXjqJ1o/YPEz2XJxr/DkEP1yl6Q6x+k2goJzOEhggQq5eh2t/pwJUnZ58sEOhHcs9038J+fb
YG3aIk2ffOe5Bnindrh0rdnSK34BnoXa5JojesMTSSA7NfcIqxCLDBtQWjHPdwisMHFCze72GP0/
6vpoS/eZOKX91MEL+7CwE0PAovc4X0i4DPz1NN49kEDRuKTfoRufYtx+Ib5/Y1kZej/kvx9nRtBm
ZE+WdvpDeU1eqBgWVY1vMwLp2Wp/4r3bjLD9yZd21Qt3Ie13aZyT52j55W2lczNV8ARzE/Emwrco
CG/J9LeSH8EcF4BVhO2ptxeBw0vGxVjGic1tdJ/8QP7V+J9qKjwVxVEeemoRfqlbUfWd1tnb74/V
zB3pArSGHCwwNTM7x52Bs6c7/KuOy0dAXOtoL/rdr4Od3PE6VBFmvzsBquA3pzEz+zjLD8xbuDHv
CapHiwq0c1gLvD7xD8H2LJNIgLE1rrC0IOhVDYbhqj2a8Ycsrt5k/5Fdf8r4p9vFgjNisc0R3MJc
X86fLDyUh4+oPCk+fkPJ+8NUMtgDjGenHTsUkeSxPZxLEJ1dY2O//qzJXVx4lACdW5AyQL2EjpBY
peT/3xLoVyABUFmVl5rF4DgfKSSLv8UDzTJgnGjaYB0OFakTMoAjBRcye5v3sei4g1uJTw8Jdfj/
EzaagHnwyhDkUVGLZvBWkQ3e5WrLD+C69yPTH9VJmzXqeoIHpVvnLlabyUqKL/TxUxx5f9brEnDw
j/V15O28GMv0eFdnUI1w99d1s9LlR+qp/i4bJ33scNtwfZdAZasjL9OJdXHMBItGfZD6YvYqgic+
1JP3N1MDsGnK22l4SsjpkBgaNB4pH91rD0bGgPGUY2jFq8RNb4GMdaqQFK4hZDR6gccDOYXUgOLR
JeKKOoB/yVpO2YjJbul6T4ImAIpdTV3a9qTyfgUY8VTMri6bri3/fMsSXaRt9Aj/j1mDqp1fQxtH
HnvdFGQduYHg/BAof4mqZWIZjkoTfXndxHpAGjof/YJ5wCl/Qq4SGF3XOZvGXgMzUAODkpX8de34
MJoqf7CPFtZLybT852VBhIr5L9oJBX4C+srTUFOTGgT4wuu2zLdeBvLNm/80qHzcAPtfKj5jI0xi
MDmMFSELL5yfhZMYA6bwqn9iTqc2c6qghKJDia86Hy9XSm+aM9uhykkJ199uG6wZkWH4CyN3tOl0
3l4UiE0iS+N4gfHNpq/CLPFZhxpyBKEXMlZT72GHIwiyUtSuIkLkFD0hDAnC+ZFnWcajr0jzyiMY
LbQp88g00FQdRdnRArUejMSqHbcNEf/A3fuyCAWJwV7/eMK4TnC76AoX7X5fNUVHq5zol5TYXjRn
aqex3BTurxpTEN+lxtdmmLpMsP951y0D1Ax/n+XyVSsS/KEwJQcDfrtqXm/Oa26bJm+DxN7Ja6/F
QQkDfILlTCAc/8bDQxaCkOE/LzvlzyNWzaAVA1HaC9PKgQguubnoQaPVXiUbhK3b3zaP39KcnyGu
8MqRNKN+XH2qO+RzcXtEmDVPdKcntT5YQ0xSFXYuuMT9C0HLZdWJB/NGy7Y9JeXLok1rnoumjFW9
iIp81EWhwYnc2umUd/dIU3PCoWnqAIlsTLRNwB1QsQmJmqQMmimqUCMT9HEyrxNN7ugsQcpMBq6P
zNdRQd+Kge3hO6nROHeexfRN8JXZPPCSf5qT4FwIs8UFwYDHK2p6pFqGixJHEihGr2cSCVipGVcZ
23O0QkqaGQjZFG/D+ct6RCzRScQMIAiHQ/Nvtq3LL8eIbPKT14jDRUz/6LdRRbSdNCy242jIgS4r
/Lh3ghnJyTLq/7Sw4sE4aA3l4fBp59/QoOP+5Wn3+WuLGCN4Qkk2wet3pgjRgE2aMl9xtra5c/Xk
Tt72y/DfaMF3TptjnNbgFsbfGHrMHnDrfESLnydnp8WK3cEnVm9dLb0vpe+lJUOHqEBpJ08e3CYq
JDmc1eigxwVS+OwPeUmN0i3aHgQ3mNg4ibOrC3pccEOvk5NWwNg7CVAiZFd0h6o3KLisgp3Pzh7c
068rDL5GwCPUcE3mqWAxkB8ts+GqbcW5d4p3FNSJ5r6FuqcDzxYwDJg1vRwkwVvL9p9mJgIthA9U
iWvdNM+OQibDB0RezcEVDio/irGQVHt8uNm3F9kyVfyZPSkXojNTmPJyZPYgHOKU3vMoQ85pkzZX
AgZeAqdu6r+83BPZxD5kx6ZyU2XqvnLd5Nc6sxE6jAUQJ0oLH3BAYifRI+pQ15mVL9VLxryAFvYo
ahHGhq7e2G2fl50RW7yuEictIRqtGczWWTcC4Yk2wroRm5UMKDnoOKmd9R7FvAal2/zrIgsCb3ac
AqiGApd5SLQxA7OWfJ/NNXncmWQaW6KYCF8B7FKfjtkB3PGLQhbPMqgdA6LlvRsYeFpyrMShRJOW
Kbxqk3QLQw2VjAHG4QCdQHkCp0XKvFRk6zc3pw/N8aOLMHFH2MOyxqmbBRxSClmb7KxTaEadEHlf
pDqOxdnEqyXcQIZh6cPdGRHlL89tVcHQ0qM72ztVq0YMooAHyEa2t2MgWgKfX8vAiQpSSiBRGXV/
qfOW/h1P81W6QbY6bIM3VvZuUFnMP49i16hbYYQcDQ1O1VzI0D6TOUrfVI4ilyGG2IWPm6w2uSAe
fiflSHnodAN1PDvyVBNTMMB1RzkrCe+uCIr2oy+7MUtM6Iae4CgolcxSOM5C3NwNnZNU5lZ1aHoQ
/Kjj+IVc0iAt5uW0G9K3g7De6RgUV6vFxWS4kVP6oJwsGTBNxQx8VRn0Dr9bSZ9O/w2glD8sC8EZ
nv/wu56RfOyU7HCH7kchH6mZInhehUvU1IP5+x72SGgBtGLcg4bb/YiIlbaci4jAE2UYfWZIgyLB
7x6vDPlHIUtrNqIIeORhQZ1+ueROQn3i3rG++tXrbOu+qLCp+9LbBCDs6tCBHhz25DW4y470DQyH
UW+I65fRLFsOULwuC1ofdkzi/bcc6dfbmkhwuqtVqSslNPfFXeMJFcN8odLAqgVSaIlQX/6cwmFt
gbuuEG3aZ/qSvS0CHWUAFwqupGI1FjXfXRQ8MhdtB3qwboozsIoRv+nitYIlFgKDIAY8ljL7EbBE
3GOX0yR9si0MBXvU5LU2GuwMc1GVmQkDI+VdUuhGkFhFyLKLcjsoWX5KtX/WXc1Fdhn3AjLwhFD9
cjHJI7H4GdERO/5xr5aFlmfbRQ0pizM8ELLjrxbM4FnMaGDA6IX3Qqy0OMW8LRAhew9C9PA5oxJq
LlqdkO7ju8lJ+oL5+tByh/jbR/6KDpaFl7600eDNcCFnw1EJ8KWWA5j+6MEDdpK3rl9DQQuRz+aI
lGXdAXQj7OXhY3XAbxB8on4lzHcL/FZFGXWr8l7OQHnnEdLMFXVZ7R33asAF2fS/2p9aEFzHWpHF
ZUoM/xlLLcrv3J1HmK4yDTVmWzyzAbPfEH92G4dKsrByen8eZyIUmLs/ifs9EKC8abKoaApmrtex
z/8gEWyoYThIyqOYAVL1iDqmKMnhltKYfOmJY/QlaCw9luU+4RAAJQN3ZqtO/vrKAKn6dwo+y8B2
m313ORLKgs8bbkzVxEWCArvLbHbUk9Bm2dlCV4S3GJxZyFLAz9QF/XFZ+3mXwkU+Zk6KwZyk1V0b
F317opq5hVW0ZgR1fdM8ke0bOwvHaHmyhMC4rB1lnQxu88sTnl1vCmocDETCXSXNjqYIyJRrQbKA
TvVH9QsUiE0AJxNn2y9gnonUQsPMWM3qr2/b5YzzLB2s5vLLoOLI5XsKIWhn0dEeChvhHnwX95QT
5Ydcj1Rv5KC4iS6C3ywOyLkSBOlnfFQw5/FIZQ71GpQMaXgG0+B0BInirnkG1RZpvTUBYbLT1uCZ
QP43/I2SRTFbOHD34IFK1uydiHbANfWgWJSab+uvYsOBlDHjYLgDZR0Okn3ktpPn7wFQI39SeaWX
nhZaN/wQMvvv2ynvpu9+Fv/RT5mygRrxjAv4n9vktq5ctjzFV9YzwoZ9Oeoghl1ejevINypkXI4t
8pt1oNtRGOsclR2+3ceAjExXrgrizkq6rvonrxvHctNm7XMhK2KKnE5EqdSrLKDyIPEFMzphd1hK
mEDU6WctBKb0htHnHxhmDeSdcfknhCZ0A+QVTqbDsF70QC7x2UzgQRWdaONd3j2oXW0urRbU61hJ
dhzJG+i4StPL/wR9O91gYP5d6z0tECnna4qbzgCPPpWCeD4qWrI76WBSmUe9HWmt1kEpKsr57a/y
Ji8kfDhwxD1dQKh7CsZ+V5MlCDrlGvq9qe1JoISH9iOZs4SbOXnBDa6P98JY/mKl2vXlRh8xyaJM
Udsl1ciD21O0FL0bnT0Nci/0oVOGUDqphPtAVSal4dQgb/xoSzhfb0+8opPKHJsd8tYofX+5p9C5
xfCylS8wTsg0ONoNC+mDpYVs2OdLxhwpqP0oj8ZlxGkMmbpl3KYFfNK233dc2rSDhQCZw/Y8+617
aAp+j6d672TcP50qbcnsY8sAtK7U8WzS2hWCmMnmBJDmnQZ3ck6nyjKBr/nKQGEXcjxMDZhZ0Wxw
JO5auGW5Yar09Z9X5f3y7jkZvXcUd39Wq3oI3al23Nny33W8lCCewrhDHKReSheKyT2SRxxvnjK0
hMdvVTXzhEYP7WYtY9SdclUtL4MQXrURIS4GoCRY2YHLz9iWt50DFj5JNIGS7NivlW4xVkZwKriA
1/h/DGfKkt2enn2ShRJuKmu6q+HosUkKqCHtNLLALF0+87DRr5BxJB6MMhMzGotvkAiyrvA3iiyt
Rn61d6PDceuL41JVCJnt/hn1bNoDdJ6QT24rBZTX4zEPucpnkhk9ylnMhpjj+8ZpAUPJ3WPQicza
+qQXkuVm/+ndtpCIqQUit+KyLjafAjNR0cmJAlhY68pQOrRpYo6M8JsSqHnLSULFoFtjWJkUOUmP
KyChyQdy1P0IFA3WxmlMuOX/J1NDr2bFSUerSteCXUS3qA4o/07s+lbR5AsuEejke5l0mDf4hHBt
nMq4Un0imKJoyCtR5/W57oD4W/lVsb3WxpGfVqYlTkigPknjQwwiJVsIhvsZqQGe8Iw2inYqShZf
Ade+vZQVi0vQeeNjyH3ZxyOGsDLM3gtL5MyJEipD5AhkOxbtAVXHNDNjzDqz2qoli6KRRkADg6WI
WJwW/q3bwFQ/1H82n7QpIDyaPoHB+RIHuGcF3Yuw52wukNkobPrwWBB86tXjrv67KyQh9OkS3TzR
QNGxhVhOSm7bs4HLSsSbh3QKGhgH8/lxK+K3Fg8dYtB6hdtENlx7fCsXoHw6caFYx54qdUScFKtc
f8Pbi5EHcAyiyc7OoashViNbYRDtLgrNLwbuRGyb0JUkxQIjkHpwUmmO2lpW6uyY1PLtRsdnV5E4
sGEiVn+1KpXNEVKWRTUMss45geKnWgbhxbK+rmRBVp+QGhcrIWX/BjZQ0UNzp4gg5Zh29MDVs2lE
B8sZdfeeaMylpM7Y6MAXCqVXUlUH6j6D1FfAOwHrSvbmtrhDFjsXQqyuj21wExl2ih20QXB0/IsJ
E+XIyKbTfcXMeT0qXgyYHV8cj/qdw3un1Mqmrjn5CERffEObxvfpu4daDb6q9R1wgsr4lUB40QX9
M31Y0o/vQI572dEklUY1uMEz1Gb1qFZN3z+mWbTYrCjpgPqVo9tybgxVMqIbWUADObebqGyl5zOH
kC7f+1/W+2Q49GlUAK3Z3TLmJzMQPe3AQjabmRUGge8RAWEjwPUJUUWMl4C3/TZIdkIg8PnSn9UB
HVEz8R9lrXxGPQIQPtK69G+VPfgBVBKFx9qFpJcmo20VQhf9pe4nSj1sHF9xH+Rpl4Gfg+ErPWH2
pxMZbUNq3NNhZj4nw/h65r2A12ahPiYpnqPOrweVDTUBkqhMWmbJGS1DwsPcixfK+JsIO1EnFy42
/eot96WZFx0624GZBj+37HTyYzPYeEG2nZm1C45znypQrRmGvlBL0Cg20mjOvWZqcDKknhoDuAYC
oRlKFr8Wbhe3Gjv0/JRVLDro0d/5FLzT9/pvzVHhwfEZ/PyjHlLrNDa1x7vrmOazF5oJFJ/I3bVF
5uwzxb43TaFsV/zlD39oFAW50sOyrQ2FzxAskO0pv4drSTt1on5vtYgIh4FIRcYA4JGbEegQj9iL
YAHaPKL+qGJ/bICKPt+AxKlPxWx19k8VS4jJ4ITZbHQx0dmDwTy2mYLSivwczas/Noszix9r0LaM
reDrkfRcHoFzfu7cdWAMRmi8Hm/5pGgH68WmGwyDEJqdK0TWAwalxxLQ6jyWLLoHTnZLw5wVisBX
NzpCiRxfZUcdrqpaosX0Vq4l9eL5J1XctNI7N00ZQg0CamghSUudl0SXTv2wk9fqkjb24JlmnC9z
w4A2iyaKdAI3kJL7UnbYdpclZNQFEGTS6Ndln040/cwKpROJs2g6rSp00Pa/RFqFO/DE3558GN62
eEIPoNl39Tb4SLvEXOAvQmeOSfYrTmcWI11WkGLSxiO7r6vArLoHocceP0STCmGw+ZrEO5Lau8a+
bLX+jABaF/7qGh27uirCqUN03mC4EaOeaLco4A2rRVMyFh6MaQqFjyjaneV8X1W5cQZHc2aZAuES
ZAMGYRTVx/EN31LgndQ1Bw/lGyRZekxQS94E+miTP8sCKf79LgJW77itpRoKKcWtB8xBPDnd2tjv
ezwH8bnmXIGIiHtmZmS7DOhZTNQlyEB072+N4QFU/geQ3nwyW4vyD2oQ34z2IMPwrhUBOCJHqSEV
DH1ZNbpCvglBh4KLq3j/0zSGByhAFY/afVxJwpnsE2zMjx5aTiyC/Y95YY2gVbma/7kvMcC+g6PK
YJgu8hkhYzEbfsQ1GGw3N0n55GmA+BMFaDxlPmVEmDbGvo9IJsvXBJMKEgCZ9QWtFW3ZWn3jJHqU
+T0WNp8x01n8nZ5t1tF0UnJVJ8oHTvC5z1cj12AURT52PnJg7pVBTOrc/lfHcBn7DJGm2BTsF2Xu
qOKR9A8PvEHrz6SBL9xRd4AV5AceSJk+cwFfKG3ZCGao07X8Fo7PYBc5KDU/QHtNX7fJh5Yz6ZNV
TguNfgYwPXGFXvicJVrTalbQLLnsFVF79iLpGb8df/3FyHs/6TRuaylN2689Rgc9QJpRX/Yu2+up
0XBZg+vVEnyV8mFz9ubbkn1I71XJuQp14dkNewVVyFqTN2XUDLO6bbc2ROKn5ix+L07CffpI78wc
NlonWVIyUAMMC6v73AYvEM99wC9JeWmSIa2/keJvT3MeflhB98PgND0bHFxANE6Ledojf4GwfJpC
2fr8lEZ4dEt+iLjbXcXqj/oZtI3v/GDibWz2KxuLJFRyeE7IYnuHRl2hFBnScmuhUgV5/3zjQ8GN
lDbsZo87Hcj6oKdQQB4Wpyh5vlAS1Bu0KMabmd4WkJkLExyxNhcS3jJ+mBBdrVmg+bT9mOW6y44H
97id9Uiy+S5sG6cUXrHRdUfe1B3/U5CB28tpJmV5UJ71m4bJLk/XihqblgxOJHRdlON40HZZz+XP
0RIDsf6vIRsP4MnhwCsenDHXZ3CNglHXG+AcaMN9t4QvTVVX1kFXnB5V8d8bCctxwT9DGIWxJHU6
U+E7aVLxQ7Evk4GQp1x9QIa4atviebp1BDL40e2YmnNi/0k5SLlHI1Cdw9EyH+nWRGnwY6LQxf63
YBnB6L7UAeBPwN7HxAWMFzIQEJbvw29Rz6M0xrrQk5FR+I9WJxvhNQ2+4R88cZE8iTY/PpW4Hjdv
q0wKEgxRKSKRWYFOCM7wIbhSNgMcAMeFmFkd2vusfa/qX0stRUp3L4oWAHOu6NeREurhHLW7RotJ
nnoQEsXOXAUfv8EN84AKxHLKLtBhvJNgcro50OPxi1C3KB5KbLpl/AYzE+d0pL9Ri8tydWfJthqE
HUZXpRD41/rFT8oWopd64iNVNKBQdvB9RuaRodkKzTSPvkJz6Y+t6yeG/jPy9tAk8MynI9l9MnlU
7dsZbBtbGf9xeqRxC1Fvhv4BLHicZ3KOiLvPa9pkikc1HCQfSjOzNLkhR4TrPuqDjZIlqzPr4+Ql
Sx4UFobzkpSRK8CKDvL20tTw1pSqEUe25lsGlfTdDzMGj5sZ/aOTMZmGihUpBn8i4+sfai7kKkhv
bGxwpitqjEAR+fOs3irovXcCHoSWQ16ONDnl5egFJjny2GN77b5kxvmzHcy0tAnvtFftF8QD1TAa
3C0H2JUyU4Zktb7JvmP6N4Ug02UEuXQzv4xD8r7OYKH5Et/WwazSU4gmhDr9RN2ZrFpUW2e8aU0A
poUgze/VbGdmWeTtx3cssUDB5H3Jj2d+0su1ZBCG5iC8+64unsBEfYflIhEZ8DRyKh2frq4vDq4k
wjECaucLjxG9S1fF2+9OawDDw3CBWAEEyTowCC9Uyn8e2c3E+biWmKOUKsLKSVvmpU5QNJWPF3bF
Dlfc45k4QCoaRh3QMbECslt/M5Oz9K2vTmNMPVguuJvLPp6CLShaUrnm7UCLSr+xfjGPlWCOAtXt
xRajDncP4HL/IFHgJYvv+g32Ckj6PKp3C1pcveFh8FFgSkf1bSaY0zSHlPJW3NeP9SEtPdWKvbYW
m9tX/LCbgzANJt7YA4nMFmgDUQ+WQTvPvpExKCmAwXbeu8DXxpAa8ze5MbLiYqcPhITnvJP0ib5q
Vu86tpT27sncgG0kqrOIsC/RE7gq5F7XNcoARqsbq3prBaG2eIqJ5HVFVoTXNIubanbWKF/gmNMD
igF4FqI01PxbPaoB3Di1HGnTRD/0+VaIJ2WDJzHSfda6PoxJR+594zEX4MgTyURleNyBN9XSDsDL
LkdqkFObvqM06c84IOLi2Bbav15QVzlwrT2vYJl72S5qrPXfpACwjPXmrPTSk7O9HQEVD6Rcjxr7
1EfJehACTMMQ4+ZOOFoxJaI8UbuT5cZkMD7X4QD3C46VVZTIXc0sXJ7EnJoKlAa5AIT5TZTMSKfy
o24MiSAUbMIw7LAftYzdG91dOG9gJkChyCX0wgz8lkeg8mGru0PgGpOCZjlRYGsH99B190/uJQXO
LcgBfGT0XJ/7KAIIXcjFcuHoeY2WiYYXYzB3tbtClMA5py2+R+HYiNnZQFBik5YYM42DO5HIIc5L
9nChcOMU1+2utYjiQVWI2ypKMV1EcZDLJZyKw2wJv4yJjT87u32Pgl4MU3MvrowLlhdrTCMGZJpJ
hVp13168XRvSmyVPlSC7ZGB6IJL/bsMUX4gynysTk9LzQ8edd4KjLuZrAGSASkoItaQnWjbRntUe
PJOLu8MxDeXFDkrJsAOoaCjQ4iwNnhLyBsaVX8AToUC4ZKjImym4W3TD2s3LQ0lAhfqXBZ8nY6Qr
BRAzqLt1/7bCzCFj/hThF5s78rrNkh1rl0KtFlnCwuCm/J6CvR/k7dgVrZa9+sYx0ZVs7kGWM+wz
5EXGf7FDqCw7zeBKfbvErX47G2YS5JvoXCXzbJpztnb7mNTJ+mbOHOdEr8WKlhbh6dt3AIZ398tr
5MCS2hBLYw0FtSnmPMIyGA84p37a1iAw6YO8g/CGMrU8iaPDtKztgjT9aAEyzyqP51wZjBSwIJFQ
iciMzDYvJBI5/LgN/px0CfsKsl5scn50c92hmn4reU2Epe6rJiNW1LtTZ63QCus/3qucbnEH5ogX
Z4i5kuFkZKgbSzxtQcy0zvDMt2ZWidaKgUIUBvwjHzs30WX3Xu8h46JfAo0OO7IkT5zJsRsA2D7U
bBixMfhqSXeRJnToI2IUndKuK4bkWpgvaDk9EG+PcMSozB08NBFqh6R8MOq2OY2OTY1nAMcP9jyw
5OMrWTxv9uhjeKK+Ve3+mhtD8QBU2tDE0TkyqIDGQwgoFl5PR9dxZDInCYxFJVEvKIA6W8j9LU1t
WWXT7tt4PGXA0+ktmaSTTh/R1Z8fCgy7bjOHE66TKRCcIw8aVwnQXPKEikasj2ohVFNS7ZYJu+0Y
+Nmk5ryDll6Ur8yTwpf2c9q1/n6eBjQkc7zA38+e7ZR228h0tZ9E/kuwZFQYXiZovL9qpT/Ta98L
9IGk1g9oc6Q8LPzbI7vSBHiaa9/b0kP87pTk5N6mYlKhHqOwPhU0O8H/MtBuLfIZnB9iaJ0ejEk7
MMuSjvFlbKPDfzNU+Nd7jDMgx0xZhq8qhGDz+qvgvI++6NJrKejRpevOk93vnCTNS/DdYkHviJUU
ccx+EjxmhU2NAdnrdotAoSt79Gd0X+prqtjCkmpOJRHUhOXBSLy0d8Bdx6BzwJTgtgOxfs/6FXkv
kqR2IO4FCYNW8BruS2zrxBKwfEygerLST59yG/mMTz3NJ8z05HPohhZ1DN0ciOrSNRHt8npklGUv
V3fr+p6ZELDZywdLmQSla9lzEhK4hCo2D0AnuZcDmhxk7qJfaT5DTp/Ibbfroif0S945x16P0uJz
uc9quRAA0khgivyzcSJXyUjlAzhAPQCcOHTB9dRw4qo14Z5gM2JOeLn5VUwedWnwqWvDFSuJNK5g
5jLqX32q54SOrd0OKb1d9qSzcsXiCZ7NRIQXXJx7aYphgnpdIbpLfCbNu/ygqmVaw565TAMUXO9R
Rj3J1kjqRRVYwa8DA9eISAmnL3Am/++V6/fmDV17bS8leEbzHenJeIlqdyVP2w4JDvzNAswwM3Xs
91ZkrAm+c1DIbiB7yJrQ7lnN0Df0DNXsvAvf8+j1z0PmoYPHvc6dJczzdVR9FvQQO277E/KbksHI
DOEYIUonF8FJ/MhyZGRpAGP/Z/0vd55qhkELeVPMcIF0IVvLW3OLf3SEs9wJZYk5gbk/ZVnL/G13
ivSHFyeBqOmcleF1hC+kxr8bSfG+PjtjXi2BDdSpq24fXPrAvV+1cPOJoP2M8EEKH64NjMrGuGXU
Mzqs9URhnpzkJul3owJkHIlDhJHwnAZ+wViEPCC5zmg9TsYXlX7rvqcsCRdhWBpL1u87bn2r+jmF
9v/Vr3nMNT671LuR7t1u11IsiVNvrYifVQML2XVQ0xL+9R7W24C9wSVzL6OBwgNn99Z1AGFLS7Hu
mQ8L44/+Rp8wQi1JZlnajiQQjZAEbWsMQV1rKdiwVgZAyEJ61AIAqcAuh6//YfR+IQh0iCCOLiA0
Rt1bHSsdTGa2eU5DdeQnxtmWlP7IkPp/xUPoiWMIkA6blZ7/3ZXstg8kkRCNlLFyKdFDX658SPEt
N3S5vTQAzzr0rEjUIPvCcPubd1ASpHRV0mPn28Sn/N+FQ+aU90TFYYbP5ooVUgUMZW/LiIuornwn
zwGsMXXySyfejcAjvRwR8dIJZMkfFzk7hq/5Gzug2Vxt0xV/8ZmDsJfnD+IaR/2VozAKK/YUXLJj
5EQWd6ppqfSOy6cJdZ6ZZJdfOpIIhzfiGcbUeyq5ej9SDmOs9+0PbKtaI+De/6aHUBxkZlG73iIm
26mUrg4PM3C9Ks5y2zuBeYsF5oxyA4+36BJ/kS58fh8xV5z+kiX+X+YhMRDRKuPC67rF5RXmEz7d
qtkD3LG6CfYpnsY32lC+UAhx3gBIMNZU82vvHYfazB8Zyn/oC5BI7lCUW10ojY26vaIm/+wmG3Gu
MTKckjG252MJlhYoMgBMVYbTHMKqTTQVMGUgymty1v8Ayy+8hYoYL3KDOYclMTsbzIO99Sp1y4c+
cqi3ZHkkzW9Vc30DSLhma591B/mKQ4XIxhsp+0AQ0Z9/PQCMlR+voog4WysEXXqfcudhApW/KKPr
PSm/KXiSdt8sR5BaQkQVqSuFRfCiGIbjL8xsEIDyreVVhQs8O7IzeIFMuoZDpbJcFw4ky0M7TA3I
RXUcN4Or2ppdN6CBwz7vsrddcYvLils1DVLQL5fUtZXgdzrG9sDwJLnjjc8k2tl8V0d6K8/4DIF5
bcykIijAgzfVt+fNu7oPIMGriQTq0mGvqykuFQYO31S797YjDxtL3ogop3P+mOeHRMYSNLcTuicZ
Pw7TcV3hNQgWpV8RfegJZk22WfB+HgCgBPXXW+xPqAJ0DmG/Ksc+h8B8J2oZurYw8Ber0ON75vT9
Ex5jN+LQFlmIcPrQHfDsgTmD2JTQUrdllyrdJqlLwa9W+uqns9qrOL61wKjlrvAJYhyDZRwgbI+z
kpbuMpZNSshrjluqnMg+A+3SNf1ALPjIRGrewPvTabRr6FySxxUui3GMgkauyQ73Czr/BNzRVEZc
foznzRgUVUjRqnl7DF7comsP50rZnC6keq2UKdrfYuSULJ3OX8qpM72OB8CYyi28Xyy7V7s9SgN9
R5xuOWJV5HEmUhDpallvzzQp5dtSRTIQcrWGeBOYHuBYFh3xZKB4SOXsf4zz7dx6DO0rbIutreIm
U7kRxxJu9VUflYX3ZCmaKliQjWgdZko+DAsHCuVXu8pyhg1TDFvAhxJvhq+uomgpcgYtXNVabr5i
xdEH+0JIsrbL41/4m1daqq5mtgyqpWo6uV6S8BqsFEFHg6a8Z56IXrAySLnvrJfjsVpwESG8U744
mpZrjyrcH4Ofp7LKE07JQxzRrXJh4fw2WAK7DzlEEOWDgCY21qodtpaa3zJVnY/Bs6efivS5egCa
pFkzM17yz5Dhp+cFWZXm1NoqE7Ar/nVGgUOMfM5YLX4x3Atz76Ht3QoqxsbOSqLkhmA9zmn7wtWA
qkIiekMwUHGoQOxvV+ob6Q3ZRK7Vv+O5lP9JKeoSMTnXkM7g5VnuEhTVfmh+RpjekNbswmxqswf1
fgS6lAeeNrCNqSeqdvuEm0sytne0V4blTIHcU267KTOYyziQPLaIsIekWK6UiccsStxDoaHDCGsM
QBrxYR4gadgWLpcHXlYurOMqcQyoB32pQMSOC3Iqjl6kMPFAaKqVZ46tbQ4lYhrZU8axS5DQYaAW
3LU4C/FwfObDXOkEeiWNq3PQw1eNu4fy+eXWsWJosTsMi0X7zwSgn1fQKOEd3jCCASqbsoSyD1wB
6Mhgxi+oKBAo4Q8Zuk9QkR7CRg0q6DMc45awj0HpANeLPg0/ISV15GoxANLq7fhukc0shmuqLRAe
r89igDVPgzsjhJIF4FihVHm/wBr/Q3yiwgAsIzfr3LRIuQ1ynKXV9MWZcwXJXEe47TAB98cSqj3z
s24LiIP5BkS3p0lPD4n/VhnFNMIxDiQWxU8v+Q8rRC3uo565Inr50+2Mj4HzTqVKZGybvrvhaHSa
pZfcb8U/vy2waHZqH7q3lmzcAM1p9kXQUyBdT0xZ+ViLBWiUMiVxpPyZVVuc7tZEECIxhEIUlko+
uYhCHpKBZGXoNvEe35vBJlZFY5bW8bRjgeVjABovTs6RQu2Szb6vLE+y54yP36jbN1QEMVlvWaxk
QH7eXFjAzNpF28C7doSDMFGAEexuunRUjFFOejCSNC1PgMM+ggnInt5Zsf9jAKoTG4ZBtyHb48l6
VfVRK8G1vqyctXVcB3kXsa3sHdU2GjWRG28tWGP497ijaUn6JbKGlNbZc1eOUE4MOcv5GXRyy4Kl
hQaEstS+uUqPRkdM4EiRSh3FlS3OqYxOCL+U5B5ng7pC57BqFlzoMAdiNj5kD9bvrgzgxMHg6YTB
DGZEVdNyNepXFhnJPZmffuyqs1zDuRWc5xaYOa92U/HQ8Es2oTDFDQgTfJBaIzOUJoHlMI0t/5MD
wOCy6SSYm+LAAU65hPFAtoG2vp+3UAMkbTRTAUFMei71gHQZvCkrR+PFP0JmrqOU8iCl0f37TwEZ
OgjJuN4zZMsl/5ICxMG8XCKjuTlDIb56ssejOZHQNlSwfBDTXKA/sY7GlF6l41vwL79P1g0r23Tn
MqjnOz+B0X5pipkLcEoyinrlCKCY3Ud2r3XGi4CM5EAm6XwiYWbON67VMBHtszp3gpTrbBWELgOB
DIcG8F375b8LKBu0+cmCRXs0zCipjb0c32Fm0DLee9A4iZJ+YbobqD8ziOAfMd2UaW33IBA5D1ZQ
14eI/UDX7/9Ui4ZrRSt54YAVAx3f2FG0kZi2HMIsozKTm4KkaSJ6muD6PVYvNOZD+TJo5O8p3yrL
VogVhIzGsf8hN77Swv9krwM7BaQ9X4bwJHAIZr9hB8eh37+LGwUuQxfMtw/levjurj6v3cuh1lAI
Axfpa8wvJp+3WzdBBQ3Arq5TRvkJZW2C6TCMMWZCJt8zHovi45R4Eq5kNu+KinZXwgYyOLLBe/u4
FKIjbbrIBMkLbCFreRrI/VlRLSEexxPKMzib+J5lfhG3xEvurnOLbZOPEvZZQ3LeRDY9nVS4re1w
mt1xi6Ry6Wc+SEuZIB9QoKkHlIzTaVHJ9Ym2Xn7ugv7fVC8yDNYTdANikvUR/Bvlfn7EY/uBgFCS
dXbaVcPmid6F48DajZ0XS8e0u4LnGJMMaBE+ChYgMWzhJM98CnVn0y08FowtgECfu5g7JMWZWYrl
1+zG9Xc9AjnxcIFO+7RrYwz167FFIGH018df2hZsGqEidLHcDHeIEL8GOgSwclQrpJzKulOK6qzj
4p2EVmsUxPeIJ5L32HMIoYC/rghTtzne/PGmW/IzqqdXEIBEGT7vrYLWx9MVgjw2ThsW/mK8SJ/u
ked7z2kdFbbS5cAYICfLVqlmiAPRZoGLhr0PieAjuRWjQ2rjv54+tG3z1jzz/EK39f8zyO8glXXR
BYq0Bf8gN3A18DaOi+foXNa6RN6v+CvTESmSG70mW3hMJE7SEd2j5kfVkmySZ2zmWGzY1eWWljHL
Hl9KyvwzEKChCGcBq9J6y5rnEgqo98eOzXRFALns7R1D7edrIRZkfRYehqBPDvFSQhoc7k0nyb9/
wAsbN7Hv+mGzpQDmDK2quwdxAizKv2rW6n3JT50qdeJEIkwtsk/FxIubvPpB2Zku6ClkWBU4J9I5
/cycr8KtZKP/ChHxruWkPjw2n+IoRCX+epFHTzKmqHMVNZXDlz4kPoljAJuYKK8tbz171/h0lyJe
VGNrY1Luy3NhSBA7kPSZt3xRtZfEbZ6TXSNEvLQ3pEoTYydlWopesTQuG6w1PqD8wcor9iwNLnuI
GL2SFCgFVHMx4MzmBZRsm/GrvPBCYRSNVR3rxnN9ZLuATFYeCXJHoGPhV6nY+0Z9zQC7ek1DT2Rv
5P4DyIaFA8gyZJZBcv/iwfwKu1b2bzgL9OdpZhjqgJv2Zu18VnY+6VPo9+YpDqaFd3mCKRuvUycH
YRMfvq0ITrL6g7916lr+NA4Y+b64PVRzMbLBQwoVOs2acJE8OrhTBj9E5reclEa65QBK9ldLS2mO
taOa2b+AtAXkFCmlXAAyJ+5EYUpk1Kk5uRhQ98L50xPjZHXtjG790RshEgoe4PhAlflOqIebgwNP
fSXJ7/1DCNE2mO4jXhSn145c7cfRYdYGDIcR/L3VaT08iXjU4F0fPInRqM14PiSYbigp+nzizsw2
lRh24ijYglhIkyI+cGDnfn4Zlu2Y3O7GiES7Zpab6L1yhkzZ1KLLehU88fsDeuV/j7oDi3kBuyo+
ZTuy52DNYeJxoJ2noAsWAmMHxpbht6qW3XZSMyPCZk6c3RlQhin7mlspz5vtdAUCgt6uQuJHSdyb
SsR6xMYCo1XC8Le5RuQthdf1GTtF37zUcXOzLIW0aPTdQfEEVCWm+tfHeHHqmNoM88S5nUbSGeam
r7LRFxfeAl7zGVqqmM4W0UxSayVXjSwQkxpvbdoOq9J+bxc56J3Px0PhZpczMB4CPWRYdBktNuJZ
3PIcqRXwtX+NNuR+AXh3NRw3eD70fzLebbcHoKCdZBFJGamMnU7atf4K8yUQGa7Sx55O1u/krfGN
krQUh3L4vxKgqXEqAfbeWSe6DXMj0SrFOLsrDdXFPjT9hf7a26t6NwC/skgmWpaJKBHcZhaEwGtb
f0EjgNtGZvC/MC5M3kDInVOkN4UqqR52lfJ6gUVfoIvhXp503xWkS8LS9S8vqrQKBCzcbMjIvEjz
VvG9wu9/yanAJSGSNF//jCFwOUx4jijv/KK31iSR1Pan9WTyAgQWz/xqq/4vOJ/myWswn8S4GMFH
kZYBbJUvidXhV6RmNqR8zy9P8G4ew36U5Uv+32VGYkfhcy7xNkg/TO3UrTyidgzxVjUFGlOa8b8i
O6sTwJKgvG3AJGgYnuYfacyJ6Susyu1O4s7QMVt4IkaueYe9nX+EkP6fxPQpJkLkD23VBszdbuiP
wdT7oE+xLuRxtCVgD6xGnlMuqsfK4WMOBoxr/kruhxRgYnblWd0aOeZ/Bl6HRQ8NZgszewVrC7pI
V5SFYfmOeonxPaFta9VdewCw/C5jCYYB+VHOAd3Y79I+XJ0F470KaeIv7qBnEHqwI7+c30yhiroL
LBuukbriAbT1Glg9tHSNiDqrhwvjXhsHV9HMED4oFpsMtcpndUp7tYzDa9PBhKBo3mzHxqr9bqlz
ZbRy3icVuAUbO9Ek5KMzWbR0Oo99NrAPMx6yI0DpL6UBviCqJvkEHHy8j/+LGHI3BOAE7U4Zj7al
yaWKd1AYzWUddVjQSlwTucED47tpZv/dBBElQAU/qPEH7vSXrPWIydfZ5Kne0SDoURgZxefxKs1C
aqvkC3ij/lA4gOKMfewXQTku7kM1AgthNYsGTa87E1Nlhfzp97iQZv2OE+5Jfgbf0k61AP16YecS
0WVYNrUraoSfN8eXpJ8GVwWHqaQXmcViJvyxl1KXl1ZxTkFN6YOLQxLOduvW2jDpoeubU+6CebLz
P3h1/6Q2HkBratEiLjla3nNqRHkPc1SyIBDNmdHMvfwBPJYAidoA7J39oOeM/2tZJYoXuJKLQUav
MYz4oFfzhXQo3OKkYuuUZDI3vS9qookTMs75hLfB7JqCsFHvxv8JYVozWu0ZsuBjKY/B9tCBewzK
Oo0LwADnxKcXFKQw3GKy3+upQl0C8Yzs4a9erhhHMALLaxfG4bJDnQV3E1zzlbbu3qXMbD5hVSlX
oE0IE8oeUVhqjt3o5yuKrB9Jo+DVcHKuFLw0p9ctlnQYHdCccSdxsc8FIk9bYYoGxLXuvYEf+fk2
WqvD3xkFuwU3kS6FLQvxOc9PLvsd5CrCXaJgIYkjmh93oLSpnj7wAujCTmF1kEEFTjjGVNSN0Mgt
8Mqr4NzwdktiLkTRBk8/fZMI2Fhk8qMIU5ZkKlwsaXXkBkraYcs2YcgpDcAlHEtuWIa8bpekbj8s
uZ5hAGfZ3wJSi/RsFmWY9k28OEPzpyu1+EBUZyu/wK25PoJLLjwCXaLlbAOsDe7AyFSbl4rbV7Td
/5kjJ/L+MT3/vO/lLK1P07AYszGbEtimg/i11Ji4Tno+B/bukpgRVtAKIcm/NRxJWY51fohj/4jL
ixC9J+fY18UG0eetFzxmBC/KSVznuNouBm/8lg1D9wtLIUjvDpJOmRvlUIbAvPlSypH2lTgJOQs/
0qtzgfMVCnifh5RLLfbS7ogp0poVIMVY0/PR2+y0YF9eo0bhrinCFX1+V2iNJqQ8cSnt4qN4S3kE
7MVryrN604lf4aARML8lyidMeurM+2zlmwpuKYEUrc7MNR+JuaSeooUeJDdRx8imRfTRC44V/bH1
vIWkWo3RQsWh+n+gK2H371Czk2w/u0KEVnA1QrykaRPTxETmPx15CrmUp1eobD+nsgmEUqpevOen
u/j15UOw5QAve2UpjpBztObzPetUdB88tLwGi0sxbfiz3iurAzMFTmS3dMXrd2DyvqGvly7qDkWI
RZWVyVJGT3byyENXZXl0Ec1P2jUZO+hsk+AVn2v+EDHZwQINGhsb6AbNOZ77bmkRZHePeWqbphZF
vO6Udb1NMHhzqolodt+ZpBX9kYvnnFtvF4sWZpMoiCdG+ZdIlnM/BECcPjy0AvAQBF8F+dRwhVC6
ixps2CHPCLEbN5f4WFYRj4rak4wWdlEuYduJFNHcIdsp9tUrX5HCmUUU5yfSrgQ7QuG6m3p2zpHH
4scwCtUtCai6Wq2edbs1efY6Ezr+fxs/FrxLPq34AE4LgfbLkjWubVMhh6Bvc3u2Oc+UyQ+wceaB
4sGiPwqChg3QKL180woY0K1G7nJJy1M8wvZ7pCOycdmCiZy8N7LokjGUAeA/RBZw8pAyqvTpnGQb
+yjPTbR0X7ejDxa3+56nuZwuKQZkBrDf+sz9yDUbhQrVtDuERGDqIogsg2Hg+NrNzPLcko9zA896
s+3ql2opSJh+qdZHjI2h6RpvdaIj1YgLM7NZslS18G4lVNxTvdgnp3dirzfxgdAsYwSCAd+MYmet
bc9j5k9Qvx1d2nRb5KV416+7I4jzxHzwWpz7J5/1Z6Q2vIXqC+k4st04dLPzOJI5Ve5jz4GmV4N5
ZBx8BWCce/Nv3tBx8bhIPbEcMJkgDn0V8zBjlGiW8z4e1jrApNCRH/tVeDkV3cxJF1dGqQ7jwXh9
zocRa4J6i138kXNq+a2Xy8DLa5I+bdqhEEzBbiFyU9TQB9V0YGsXHVnHyYza1YDPdOSLoUVth/9A
VQZOFO4JYTippH4SuxtdMSFQ1ll2RtlNTl7aRuK+OO5KzGkHhtGdjX7IgMnoD7VOZNpJk8wl5g6S
LyKG3A6DfEhDwbG8SGhsDH54N1JcYBCxGmLKWeAntZ9CZJzlqSGuTxFEsnPYQC+IN7PQIYNZ8PoV
FIJjRb7ooWpUqJnedlQlUcRggQOrl128a5+OffomGK3vrRlO43jcxmD1Q/CKWcTlyWoUiSCY1smw
ivby74Cjp0sofflHe3zzjDCZmCEKIwyx6NI5neO+Yt4Cwg+HtOcL/hP9P7CAbjii3QTaCBpptUFR
pyzHdcv/I+b0jI4IzrLQmNqGWFS7esGXRU7WTe9G1AQ2yUx8hw39K3SIYLaAUt2yjFm209tIH2f0
eYGU1kw62c+ul8CluNefN5zHFQpIRo0vJLdPziOg3xwYENnKuedBWSCnYnjbM41AcejTJaPRYN0h
qLGiQnlYnlrAb/bfczANIt4clq1EgvR8o+/bOx8d/XNJDXyyGetWd+Uq8P5RX06tlT0MdyYBy73S
NzjdFQcbYgEsWrdCd00Otzmt/qEPfxGCc/ZslaQhvrXQXnc2TLmXEYHk6Hi0047FxqC9ykWtQF9i
TLkwqG4admjZMJ3C9VC/hNkKMWrBwNhBev6HXotREg9rZ2mQE9DEmkrHhsMDYK0I+Ij/Bc5dUmYU
k8kExjatkpyYzNKOjZTI0osH+CKyfu8zCDTLHCgNlpm6qzLbpC03mRr6oEimXKUckCYs1f2vxPEa
01eTWUzfoCPGtfihnbAh49D6sP2wWpA+u4s0xLYzqc0jiq4iG2QAAYoBDZKcLw9iouO0ENJCmgdt
pU4LXWjW21tC8tD/I1j0pCWp7VNe7qnBI6WGBt7ITVSI55N4QtM7ZeAhdnQtrPyPnKxUeuTzG0Jr
1j6NybGy0CCHInOU0G0TbKKkTUpM6AkFfji3YREkuNnqFtvl3/eJVvNTBJSEHQ2db0WzyEz8JsAQ
zvLabz68rPSM6p9K6MbVZVE4rNBU68TIdZKx1BH4jrFM9XN1c2QM5+qHumulMsX60BkmFGEfeQ4+
khxMJneeRQtCdxVifdVAAcpxE6Hz2TukT+xtfCvNzamqvfSxmJLc2MwvCLx7cmB9Xo7UJTOj8fiy
UHYW5M4B/zEPOb/RnFUkxboW4zGRT5Hmk4fmzyDU/brOJjT1PbRcruocs+wsuivbxV7TDCz2pIu6
KysgbPzw/rnoKcq03t39+WHNO1uKHjh1fBLtbmaFKTlIKWx4JNJJZbNbQnyAF643ZmzTgZzWocti
r2vuV98RyldJlKqWFMCJIiFZSIO94XzJNDfk0i0VRTD57reLIGKYs/ITT+jn6cKXY9bkoFQ14MVG
DSa2bfkRdk7YVTuydBCCB1CqooVaL39VGxRpGyCavDQuVOM0lIgzgQdhxePP2/pOUf3AfAPY2wkC
DlYaxEOt62zG849Bdepi/upDquZdiLBWosi0xTItVuX480yj6WteHqUwONpVS4uDY0fDrW8kkcj1
cDkwbaB7GJy4cb/D1Z5TJZy/k871Yate6ovS6HK5ENJ2gU/77uWMkuNU91G6x4iQiecGRUbzmmG5
N6EYdCw8QFZbdlKvZpo4fLJkdk0wI04LyXC2c3zl7PVxhQUEt0Mzuu4gGnFsCcLug/V3aQIDuaCd
b2yLPYa+X/cvcHoEU8mvvQ3Pyivl4/6nBP9vyB3Pr/Yf9WdUlCHXAAp/2+48cIQa+LhA12KxhPKm
Q9fSTTME1c3IpOxMHyrOgN2f7YajDW6f6OClc7vkL++vqQO7jNzA6MTlZE+KkJhWnvZ9ckDzYDZU
EpLfnbcTG1tN6SH+0ZJvACtD5uIznmHKF97wegq+yv4+x8SwvsHJqdpRf/ODFd1U9mdF/7ptYEun
4ilsflzVTUNwK5xRfrwdGUiBCpRlnxllxeQw0i/Cqzb2DGazo3HHOEkNtnGpvKEIJp1nU6GOko9R
+k99y0q8ctmIul8ats6MvGy4b/9f/D4xzfv2MHYaBBHbLjZGfU2FAeUksPew+wkXzsy638BALu6j
rSL4/s9NQZXopXQCnAqU6/kWSBbZX+6j28GA03806CEL4Cw/B24X0udrnuUcE0D4BqFB+vvCyWYz
7pr8L7PaK0+qDuCFub28XO6aBY2Oc+fR55WnxFLrB7nf2/bwHg1d+OpdvFXvPC3rHv7/3qVOk5wt
Ram+q9iZZD0Wza9fi+UwRSo0J7c4wGo2gWkxyt7DErejsX4cBDDftJTuEgKvlLu3B/1CcAByy2cs
vUFAoJWYb5Jgw9gLpHRTIRuOgfEzrvJiiduUwHSWDDNBkESXtVpr3gVA0LQBo9uKmZ4yvX8c8Zay
FASWrxKCFG+Ozv/Yy2Aeh8Ti8PDq4IaWRR3FwcSLHMpBU1/evlM/ok3dyxa5hQz79plA1xutc52w
pNqaTBleWYIMR5A/Fsg9daU+inZE0+VNCDWVdgEEIy+pb67WY+bCgFTLtz/E2HGE4yikT55CpCaK
zCc3kDohHFwCfrZRJnL3aUHbeceAdGjumIKNWpX8CizJn0TptjC7Jvz2Yh4nCkOHVl0xl8AQckq2
MGoluJixnJygmjYCvxGe3jM9GozrWVCTVeusNdkjfSkcbcQxMfaJNvgVrH7NPeFVdbTYIAfKRJaJ
vMpjwN20g+pyGUonEGS2UcJYy7jIRnmrt9oZ+IIW1gapsdEU7eZMTtPVFFBa8/MOucQlaeACp8SK
g8g/B2VFKH5rzxbc6a1OPYHfxjvwUXwmbfcU9qVg2zSM8DxUFarlJx+v/kYU7otJXbYpER1dOhIq
b9ReDRypPPAsehFC0thVe/I6D5s4cbCdKMZfc3VHxZdZ58nDvUenSo2Eo5CizvsvPrpZa/0B5Cny
4u4yzVUYLv6z0vDl/v3FOGGuNpLcdzNiR5BT5H9OVTWO1XUDItXPlyRjZnaGt4eOpq4qwn2QY0ES
kAqXEA5VpK1ry+GOmyfHLpunpOSEcoKJJECiycih9SIGdb/MfYyoN3UMYv+D8KPmY2cGk+Mn5lX9
Y4JayIv4Kf4oQjarGrH34wnF5aX2UqhQPACDJ3vxga6kZ0D6WjotwW3KFkAtKYpJFUkxF1TSyZMz
KWBbxy671g5ofHwYY6hIq2Ne8krwnzpjcj4nDfjPVCau9RvcDhp21WVBiNuKkY4SmiW1c3mce2iG
Z1n5tQqBDdr1sX+Ibbx1wXb2O8g2IsudeVYJ4G0pQQhHPOc838o/Tb+wi3ghEj+5DufZMZ7J2sQQ
nJ+9LOIjDeCAvBKs72vDl7+HKpBKtB4Tc0C1MBZ22pa/WzNeYvwAoWIuoRHMPUWXN2nuOXUgTvIe
53gvKCkTyhGCFBvR6NgvKUImlQOUUz+yWuq/AanZuwKyEhkK1SM+r3e2on+AgMvOp/8zrMlJUCkW
LFcl+m4jD36vV4fDSVanTJ1jkWe7wES2azCSyPv2F8LFd7H/TCV9ImXwspdD0RaVoC81UGbOxU4q
/GB32TsJUDHhM+RWl3veNHiuwg8u46s3wfD8dTJNSutZTNy2MWXZMm7FvfXYfK50ivHuy/vFuOwV
/iJ5nC8zcjGkOXZek7A2eg1x95kyCsonWcBboqDvwN10xlbX8KanyqVBW9ylwT00yesr+LzsJp/6
mKvO67pR7bJpkeU3JQ8PQq/37XmU40aiqILR0uAJbeJAAMQIuXPp5FwOVcuOFMum5oQVC9/WJ+S4
5SDUSc+vRL6rHyMsrTfusCISuXLcT5pU4AoT8azqqnajMEB83lGmvCfkFs+qxoNA8GQxj7rARggf
iTwLgSQo0XeAJUaQC3+iKimxBl8Z59CoDKUvXflkAui4JIBtrvq09hHDYXVZFG2gic+0B3BZrQEU
GabV7RFFcJuFi2g0vUuZTYH5k03zUoMJrUq/3kt4HQW8mdNwgJMCaaBLnZnqGnS2SwsC4Lhcy7TO
s6psfb09URRjZZQ8yVdx6L0uD8a+2EhJq3lEK7zCd7vPUfn4PuVo6aUuSYscMLfmBgiFZCzw17mv
W54TExvL5/KEnbShiso+bE7DDFywmQ54SZTYp/Q3rt6htAez1ECpm8u4DghBQweQHI6dIZUyB16E
3/ms3RW8CAbnm9EmR5fz91rn8GMplA4w3K4VWie2Prk+dlBjwYSIpdG5ToeS31eydJ/3yZL1Q2Fx
Mb14Duab7BQzduMuwyctzZojxuF6fJK9biFZzlyVYLX0LfNWtWkKKIah6NXfgO/Sh2k5McWtTs+/
1ZjKjH2J2HjF9XbuY1SC11Meeevgg/FyteFqtzryXe1CrDqLkR0RPYvlUDYZugRRurbOYxbUMnNC
HvBVVHz4DUfqj9AVVT1cZ2mdZDe9Kmtylm1lWMyHbGgFo5YqXpr3CAA/JJP1q55UfvE6N0nVzmiK
iIzDy6cudTWeW1lPunUOVzbkVh9tSEgj9N+SGj74+34NNS652JOUZlSTCMt+lxMbsW+FO1GM+4tu
xNu8VOpjtmXPtBH8l4+y4tJipuhbQ2WGLtVtrjKvhxTBwK1dk/2nq35DEorDCg+Yqf8t9XPTZr5U
1Ovf4ybzOPqDIIPY+2JThUPef1CuK7lKPA7CE5mIA/IAjE8PwLPm1J8TZoSEog3QIF3M5CQcgtsm
TURKVMo22V9JN9QCTXsRlt43CZtnDqm8iXrY7pI+4pyOSuLrLqgQ5/EQkhZrn16yA3Vnm5ObEmDE
BYJf/H9excbxWWdsnt2DLJrPzlr4zW4YsEsO1bsvotYiOkMntd++S7l16ealPayF93/XzvlE3Knv
SMbfuUtrfxw6idbDlYoh1LWFK9zNbpljxfSSfGKi+JDE2D9+iUplu4KBNq67yeqaX+/YmjUiUjWA
1Bh0sP5nWMoKpoPjhsIenD2hc88hKd7dH03AruPlid8IZe+MgXRoG8R1Ya6CZbj7KAi+aKSoftQU
JU//pR71Ec3DKK7xPQj36N+viWhfrqs/KTO2n20g9wkkwYsI7Jsr3ryTuhByD8w9T7XgzPLDX0Is
NWXVmeksNwjk9encQztAsoWRojz3DInOMfH/V1M51vQ8XJBpCvAdYs4mK0RzZ01KVRy+7vUOdlpE
WxS9Peut0Bbcj1Dc6F8gxvmOYz8aVlQO8Q852f6ESu3V2CVS4GpuyN7yhQbb9vUGzaWpRifs94/9
d4D7xhx4yrnCcy8vha7Jy4VMsXSsvMIIchky4r+f3JLhrKMpw4v72RJeS2CKrz643FOuAbD4C+/N
mNcdGCllyXJ/0N9NUbBleBmApcRWnsuYaQk0JBie7S3OC+qcyxsxzEckSq8DuP/5E0kYPUFftGD8
c4cw4Tjw5IZxfF+Q7aEMfeVGVG8Q1c/uWo1/pj8Yb+AODtvQ5vb3roNKXbhLpmLddfLRr2pSz5eM
31Rt2WCRvbyufHeBOSzeyAtR+W0fohjBeSnkc/L+KxanDGidvdBAWpKGG6Q6L7/0pa5C9qj9JjiI
h0ltXCMUdgGsx+KfQNFOmrLMKrdWIoOtoBndeg2LpZJhd+cICPD671Aq8yqVP0WH0sObz4Ykf3mO
dq2fRS6wa0kbwix2UrcqB9iqmeuH9iPxge7oHNMpytaa76OyiSVgV95VBjfMmfa5n1YB2Z999rJR
NUppg+do+RO+Ww0XmQc6nZQ91HjqOOmqGR/hoWKcrM0kcAopBJuhSX8f9VyQ0vz8TzW1wR5OFqbV
8xEiwdHPz9gohXIoOzCFuZ9k2jGVMdszjvX503yRSBo5LagE/gucHTKOWN4XlXn0vy5TZ/FFIWLd
iMvoiPPW4JLX6u3TAH3I/xfo/9Oo1jGrTCTbzBC0SUVb5wMAJrGYEikNhuC4TVTGy3W4pJhJGr/i
4I7acvOjuVI3kDurBpmU+OLQVhQybGM8DVi74nBsAxKjvuqdI0RkEZeaOVId1o31p48pgZN7NqZY
jnJ8RYtrX1u1wQmL9Gxo4nmNW/Tl8cT0yPUvyl18sxN3daG6ErBemhk0ldHl/CM7ECmJk9GK1aGH
P5p32XdiOTmIj68rZxfnLMyRnUcH/d++qWolSvdYa+oFVgDfr9RJCXeQP8BRlQBWbjvXo7/UW8Ry
E9Nn+KFxVyeOJvw1XApqMW1AK+IsRQ5LjjYezat8YImUJOq3Y0cnxAh2jZaXCvAZ8sZVWllpY2wJ
vSF1ZYZQWRJaNWKAYqOIZv4dAZGJW/X8ueHAl/00CAh3UhgB3gZ8uQVoxrmdrhxH1u4708ipT8h+
EqLOGQndvA0OD3+qwD82bVK8tu56YAkVyTyBp+lfEsjY0tqNsORqc4nRlCSI9vlN57al4MlW78qu
SMrl3DE7V8JP4Bd1SFKjQ5JnN6E38qnlL21b4HlN94c5zQIZUodsBmmoT+nKm9OBZrVCwrzCabfZ
m1anU7YqWpNYadzobyxuBwbpETkjzS0EI83Jhbu8NpH+x3puQaHWIqyKx64rOeF5aBWqUH3GCWl0
Cfzq5gwtcX4xPmVcMYMRWlFyRY0ZNrg+A90bONroCRrXgf7jsXXe/EwV3RGnC8xYuB2jnArblR3f
GxBJfcwpkjw3/lJpXxgsfQE5kKXhoJE6nNPUQr/+vHXrtoimOP+YtAOM+1IQOXcRZa0UKLe8q2HI
1thZz+yqIuzov5CCDJ1tmL/ZfQ6ntUVOIkEXcHsbGOhCOHa0Jj5qY+aEexlGPOReRf56WPEzpftV
lJ7HXf6igonfVY0sTY27s9L4XEUjiFHaY8EpMFxFMnMnYBvJ1IW+1lqJNpUHwbZcT+zOLK1mPA+X
3dPeudGIzKf/EF9uEoYHlhxsHvLnLM7+qIojSn2zo0wpRHErw/v76IIo2aBupduRNOAa+NY813xY
b/jhlikOjb3U9eEa4F51wewsUm3Vfk+1IO0u2PY3rsfL4gcIb3f/HQifdTSt6tdmze/9JihiVoba
JwEYYp+LXh5oJh7oPgNeiXPTerqpr7VOCFLgKI7T5Up2euzpJynKw97wI0oeA+zR+8UuwrFJ1imf
VpdB8cCKWrYu2xmTBdM3WsjfOYyb0eGrqf0iuxYPDMzdxPc/IL6/c50TpAT8pMt53Hhfo8INpaBK
yqLr2PPpJAU3Dcp3UNjE1kR/ymHI0Hcc04GiO9gxGINmvKoh0MWBPNZcXcfCOWiMQLgGlNi7ThJA
O6fXobaldrkOTBv+Xazxjz8HziNqdoXGHrYcqv+EmPtIh58aiTM++iXl8d0VwbPCYo3qa2e6UnKQ
kzwwOfDI04imGTAT+60v/yAueE/hPkrjl9l93ehTpDTxmRYclgnYPM9keGD4fk/xDxVBaKvJc3tn
0i9Sundn9RpdpiGqqeQvbG3va50TJjsyGi1j4u07Rf6v0PzdDocqA0kRf+p+SZnjytOzCfAI6Log
XHKXXgpuvPFOYa0OhJdC/28DuIGA/T8culL8EXPwpOWw/qbqu76cSawPQ3bH9g33U1n1Wfg3RXkM
j8mXd3D4ZvrblNU5L4FObf+Shq2qhvMFdNegLBh18tPRebCulZP8a4nkmwb/m7uKKZXxITa+WfFU
RTKB+OUy4MfxMfGEfXUW/s6ZMBIv2QmmUM2dGlvzR3o3WG+bJuLgDDcJwspcn8UGZogCI9O2/3T+
SpHAjA62twpKYYrHpcrrTePtxEVdSnfeIvLuBlu2LlVwkTGuBQe4ThC2jFF3uG7P78OHoEE/39bd
GKeWvi0QI9HWAf9Wz5JeE0r2qZf0C7mgtgXKPANGFmnJgc01tc3znHA+rAr7jY2Ajywea3iBDhWe
Y4+pHTFYEY+yKlzd4toWgac3H33xkl4GmTRJii2DBTsf+6uQRFvDT7uJu9vWMXe3XOcQ/RLKzPyc
wsOgw957VNcFfkWJn2H+DYf4ADJhBL9vih4i9Z4wSqY7w/Fl6zSfyKUOuW7VYtGHsaudt9Zhmna8
Z1+hjWGVwWlfCpJSRyjBRFr+8UoNzyRnULZ4ziNXNch37ol1YUMMetAS+lFFsbDNPTZYslzWBJgO
s380KJ2WB9jTsR7IYj+Uut+XiirwCT32pyqXjHkCeVOB2wd6+u5vFj9kR2id/AjBGg6zVpwyQBSz
niasYQsAftxbCGjBa23/8nEpB+A5waGlN0tA7SEg6R5qFsj4IChBZ52MZdhZbMpwuvQn8im5luiH
Zb1AsPrErDyZnRmSL1v6UwKzi2nZV5WOp+wQmBqdz+JjgLB0Bpaqv4bpSek2ROajdkKRYtUd5R4i
b9qlHZFEbjR8vm1icOHITpAM2rX3XmFqE/MzDsrX7ANruKGO5nowcWtgt6uc7BAwWUN2ePkmde9f
8Wrv4vzCoJuZbKWHAiyjcKPfEgxiNaOvcyMcwi5Nu75u6QqZikLz2Lz3QctunszE+fG5MFILIClf
Mg9w/ereLQAMcNoxkjowuioKA3i76azgRrKEl3yDOIR6y0hNEwxBF8cfDyXzRIVx4egyVWO+B8G/
14AZrA5Q1JApzO6oaPTMyNLpY8uNCBXTwpxI4EfjA/wqxYljb8FAbEfU2LuYOERIDpRDdXKercpn
wvX+dTz5Q19bbtJBLpWTVSdRa/tptLIfAfjKSfQoFZXBbZDwUtCuul9mOET/HcIq1DwmTqgc8MbL
u/hDg9rYKrsANKvquglLiUNRcsq1pFgv1oesXwtX13uyqPuXbZVZWCVF7UXgHGuJpZoupd00hwSk
eKQGbTfRa7p8yhwqGUMdG1d0TGBl4MDouKS3A9oBMPzk8s8BuRWNzZjP+GeTD99hnU2ZPbhCz244
6h/r97T/lrJQzl+y4UxwfFqryW63SI/HA2BvtCKLYKfkIVFXxVRf2AXzik9byOzoLYOI/8BUnd1x
69Lm/WfQL+6tl4GhzoPioq7xEKFNwu90Uv37zGOHmP9cAtGvjJuELqOCf1G1cb/xcBmHgJu7LAi5
dTuMH3tUAnlp7/95FPTEzjQrrsFt2mpKmPiD/0AYx2ER8Rel48/h4DJPLpI9ZX186/x51dZErK3g
pCV7fY1Jw8ynAgwXX5hCHSm/idwDG6uqSsM9uUW0cqD/Oxncc8ssPpScmw+Dbr+3lbi8omvbJDkW
g2m8a43T2v+nLTtuw2DX2IaSaSLL8B1FmfMCyPovkqLGwroxgtbb55lB5SI9IbaHFO9nnPUP+Hlo
yJf3tAW620cdV6mL8eFSg9qb42Pmcs5Daia2wGEAKGAT9LI09wHc3AC/RB5qU9eHPVlj2w7WTDBv
PA9/9Y81ncMoB8x+/WIGd/hpcpbTkYu8Jp7S+FBYOIetxgKSXrWVz5ejOpojNxIlhn2j8hfO6o/7
s8TJQf9zRp0SD4TdtfUo/EMF0sBcaD/A4huCd6XCFbWVOTca+URSlY0W7tbaeFkSt5fmlkxZ3BH/
TOfnfGGqI4f0bJ63Bzo+DYvmRdwRkiwYtCebjwnqFIAs/gI1whC83jkVzfFGvDwLOc90nM08OsPp
b10MzHJ2ZFF7kSkvr0ekgHbm0dKAqeUlXycXJZ1bQF+kLKWcjzd0GyJf/7sv/EKo0J4o9+qsEQD2
sdIlIVrKeWcYE75xpYFZ2wECieSEqZwOm4tyiLKL+Xlz6cpy4OxutX9CQ5JueQeDI+E3oG34kd+t
rxTLL5o4SZMmTgM2qsFbDnhCUuq2rEn6QxH1RAlOSyeJsIqb0m3FXhQ/S3qVcF1TiAi/iQ5VMF8k
uteBdymTJmfOwM1UbUfQoKmdgRtHfvh2+YKH1So4KE7+nU9DdDbYIRn8TGqbTQ4TH5E+3SX9uRir
SoE8zVmBAocvIm6/JaAZUp98JpKtBJfEHKUGr9AIZfHCETCirvU4O6j1Hkwd4p6bX5YaiDCyfQ8i
snAV4e+m+GmaBNn12aNhD6ra7LiZrzEvKRpYGHfnk/Ro7LRLmSgbWEqRWYgfwi5Ay2ySq/QBFxva
pyPDPem31dpEK1n6EIcrWj31cNKk5oCdhvOd6Ut64aWwJONar1SQ3weO9VElyWaE86LKNK178qs7
hOrLQ9bhdNw0CZIqgu/HZugaYgHluwC1Gx+COkdTkUkB4ZrJmAeOO7KXUa49OgxZy4O5xV/UGbMD
80oiY3/98n/QZcPtT6BAfGnO2aCrW4CaB4LksQTBAarUJD0QPN/Zt9Sc4BO3l4LGEo0/wlek8IaA
B56+S65ixmfCZ/ieGJUjOvqLZujQp8Ze3SIIN3biJjKyxQcObkhbNC/vXKOlPg+pHym6fiAM79F1
8MfRpQNQah1Q93tYLlYwI3cpLsL4EKQKAVTo/FDFugxTqcG0Xgz+0cBUyYfNFELbSS+dqdqXvGf4
cw2ZL+vQJ6PJcfWIt2h+pVkwPFWYScN/at++LuMz25wTfV3rNEZqx7h2eu5HAYYQbrcC5vA/X/Ve
Nc4mIbb+judWtYhcSup456nf74+jUPW2CSVxXAIxverIgkI53772kb7sGyH8ZGc+lG9tP2qp0s0B
CzxhSEa7N45a8J0OY+APjsZcTGbROQcNOf/eHzb5v/8Ca0ItTplGC9Bq19gJb0N4EGFNLMZypUe4
gSfnX9OvcyJ2j4ZKH5r3fnns8ZsbjMBmUHi+1FjpcaiXnRP3xw6o+AVJxf6Fpxyl7JE11NV1h2s6
RW6P3sT2GoKhIAXQL3F8j8dQLASeT+lASdRZlZAm6sB9v5rS/tZaZUsQ3B/w20AJ0DgVrANv8Aga
3vNkyJwhNb49IAqmHmzCtuxHB8iMokTt1bNv6d9a2UUf18lOgyWF3H8w65Z1njoJkW2cpZuOdF5n
TVeI4+0nrDxDheX3+DViSUwdYsbp0jbtMkA2OTQmKug+DPLI0whgmebMlePOVgplBLlXhigCkX3T
vXr5C8moRq5Cr8XhNorid19+uFF4nZB3IkE2ztYaAtpW7nJ71IicX+6usQSP300Qaf+cMRUzmI1J
9V//iQVh4yVJj3Jkd51138c6Es7FVGeHBUbnF2MhOIS7af+vCw/RPLfgTC/zWsi+u9pwbB0wD/+t
02VfvriuM3EeaOqgfwq0K4weGJdD5O04emoFbCmbLjOgcOCjJlWBZUgkC/AIpEkzN0bzZW3Ix49j
FB+X7QkQ/Cq+7lsvbbk5CymIQ96h/5czZqVx8+HRWj9ip0QbmTPh5oXQlA3GDJd59s5WcpPIy8ue
xnPd6h82MDZlm4CMHhC/Lg3me5t8DbxL0O1NSp4yS+pfcDAbZo1hsgW1EPtVpJAImWnQQY7OGtQF
bjdGJc9AMrxfdvy60gzGv5ROwLsvlHBjOixrqksKOcbbzZblRoJXzaUWNw+0S64jTrkLpa6GkO0o
o+xoU5j5khbjdpZP9kwHEpg7RfQTA9AStR4xPkRxD6FHfsQiWkG6E+lRCu0B/mHugzxAUdXIsOqP
ZT9zUDKWvVWSCnXYUv+4Jh2Ma/c2HlAJtarj1ko1fRCQl/yo60iik0ZNQJ27WufCJjSKcnV9/kgg
CN3i7drwEHGGySxMhSXKziBLSaHdWbhIb5PpUmkixUM/RZByTKrfbbvepAqTJNGEiEydqTqvMJns
L707kgMCntod/S6hjAWF4gK5oXzmja3JQunEGW7+TOJWq/MVrCtzWSKpnrCXgv8mhSkchogfGGWv
CLZOLbDXV19bLb1Tr5Nu5+/vpQBTpXM03G43/uAILQh2qjZCiE1Z7dnP72ww6ctvmxIKpJ9CUQM8
UbIuRsDLrIwzWwXPS/9roAc/VI/MQioH3usVXcYSdyvCVo4b/yMNg1qJvJ8yKYXz/53JiT3xFk4g
lmHg/xGfCPaovF7cS+eJ9rPwSSxVQWbHI8Ken5mHs/0v5Bi2qcCICcvNU3maGhe7T4FKBLmQ2Tu1
+ET4sbwdpw6tx6jQPC9dEkqN/semnJNb5tjR3bOmei0VfJ0R0bpaxyTRI2vqTQC+XaiAOWvbv/R9
ArsHjH7prc2GzmoejhzrH2CXOf9ZJf96iebQpfHDnThypuoyk+z+6yB24V5k+ZK82RpeN8N4nxTU
k5wqAUV7FX/oLOIDc+yKakF/eWpzYdSYnlRq+Ak2QcsPyvszZSoWF6kEveLwa1uqAAucmLKzuvuK
wXG4y6pEHohnN4A22qs9VaDjjEy7bk7S2sHr/jDbR7e2BBoCEXW2UZpjVZxeGuG5gqx4dm7cyLCd
2EfCVZp1f6SUjj0D2JsIxL7gOyLP0g09oxGXRRDDRLa+CUqdRVZfjNQP4v+iaFD09wR8Yn/By3EL
N4NwxCVqbtKF8kgSeI0GV3yDbRnwk4alUd3E06CaE7uHxkCesbZ5OZfgVdaaEh0n/up3lNjo2+cX
YHrK0YjxKK/w3AsK+E0b6oVVT41rma2FiEWh/X4ILUv0GZVHznQ7MG6BSoXuSqiZqgYTsaltneV7
htHkUYP5NKwKgNjMdIHl6PqnaYYFQMQsqnuJa7dRFZEShDuqs0j0ZA5U5hKfmSJsyD77xuxPWALj
VZqZ48M/QvDXoeVp2XwTkiuMRoc/hlB5obBq1ClapWXxxi4pvtU32kmLR3Tbm2ozceG2/o3tArGe
CE2l25B4K6aIa6gImfH6UI3KhS/a6a+r4uoTJc8F9269xchz5EuqTguBMCHg1DbsVrA2Hd1q3g/h
3Iiy1ZabHmF3YxeERbbi52p6v1V1mXFnQU9SHg0OeuvAGFAMnwm4n+axO1kz7q7G3LNkYScGBvfE
mAwmu44ZFSIf8Q2suTzVviqGMi9MiVMEI6/+aCcdB8L4HxvYHkeJwp1kRRWy4iKTDbC3xpJ8i29W
6tdqYt2F+sgNzu4pPytZtmVwU6qzxMDepRBZOCqhyA7okb3+M4KvDi/oL6I7vDwPjLvDPA6KnUFu
DzM9tdmy0UG9FFb4AlEprCpmCXpkKohT5eHwbutvQAdFhT5gJIrLOHo6qiKowfspRO/IO4dOMXeJ
BNGulDCKOnU0225sqmIj52yrDfr/3sL+yl7tkOB5zbsabejOTvT6ZPKSYgLeQSeQUp3Ynd2QziUU
ozOmer8zKMF2Rk++uWA1Musxu1D8UPtVPBLDapay2ISyxilSkNh6Jy9rTFMhfFkDIrLquH25YTds
AEnNnnbOWNSD3/Q1Dv+29Ie8olBY2MruSaxrEXNt8DOArW1ljv4PIRxRoHoJwXPaPXaXUmWn5HZI
+h8gnETEx9+P6dFPYYqcr1sl6LNxN1Y2U7Y7ZX5s7ZL5mBrycKyS7PQyWHwD1pQT6GH8SWZ1hhuy
LZTJ7Zxh21iMTRPjV9KhtZVlbuWQkST8x+7vg/UTPPf1j8G9PxCNOasrW9uO4lGktqG5IpkMr10p
dW4c/jD8L+19OGeu5qlwMJBGfViJ2N65+i4LL07YL9NIqfZQWIEHLnRQUSsSfcwJveWzZ0jybJep
pMIboWrJ7e692xdivJVKTquOcAUPhSHQywX3bX9XYL0hD1De+YIVHn8F1YblsgvOENTKI9jwC9z6
CKH0mqCLVaXR7Wov4xnytggttDOHsFf3OWCPrg0NSlKcH22hFoPqaz7xzvaxfo700t5YSATrfSIO
jOKTnXiDSc+VRgLhSVP2f2BT46ayxbkzLSV70kbvRMqxuR/CI7ypb70F5OnHyGpko4s+mYjBAzmy
+C2i8d7QSEgO38TZaoq+dBp2IaToZ3drSQAVlwehSlXoUfzawIEaUk/Ze9Nu9yNC2aC7qKIm32+r
cc08lRRGAblZmhNUaHgV/Hdh5V/ryWG6QyyoPVQrf6Q+81s15LV+P2REDEWiBehLWWmkMXUjEU8h
ubV1Tq5ettBBgF36fTu539nEok0oCMOZGqPg2wo961aNEdVDm2SAx9tGASVSmVK3PtWaO67Fij4Z
QVmg9BANHgivzRX8u99gKf9OEXA/5Y5H7qgJbfifQggUJz4cxGYYwbvr8EHASFbGXlGOEUbd+V4G
rEO9UcEMTRwuxcmbzsq3AGzE5Sd5H6OFUcBXPkP4PSKyrWGEiW04vWt/htr3AK4Sk/xvS4QTyBD1
JWP5LZYPgN5KcabwV00w3bcMO7zJkn+Mzm5/uZ+BK6v/LFWL2LQ2akmczYyOFQNyo8QPbQtm0cnS
odGpjx7T1SJ1wF4K/Xh6aWj4QM7y3LrX29KgH9MjK0G90L8S/E9nFc/Hq/PnpEgBCpMaIp8vTsFY
trHe8bdw7s2kreGyTlb4InZqRHB+gBqPW8Pf9THcppRVFj3COSYX1ol4SoPUJIwaR7OvJUIu08Ra
++ICLJlNH/WWXoCl+bBYYdBhpYv6dJr9cOlt2e6zLWI58vmxWfC7vC4xJeq8tGZ5AWp8AQP5Jq/9
DPK53xRyBCQZTAJT/Nd4/hVsg4v8qr5TE2F5JcfZbZJf78MeCdKvrnxzPG516fr6sZzIrM0uaG9r
sDgxiOziClWIF7RBo1omrOSYcLGvYHquXAiBWUSnlmVLIlgesX0GPKepqXC17sK6kM1nFMS70fDj
J3KHRI5Itir1+07ZLtjq84euZjYM8egpfdgecG1LJps5xrlyrP8f9R67DkpynAO9cLbuPU88k5pf
L7/3bbW4s1+CPUQu0ZrzIYCHoR6Rt5Om3aX9n5wzumy4YWDcqoSj59yAp0mt0kIw+UFkC7fzG2WG
Q1gjZbhqjer6m9ztQ7twnYH6WQkps90oi/InvTDPByFApGdT5q/oZqcT3kIXQ1Sk1xgqipt0lZbp
o3bqMDkEG4ZRp63IvLafipVAmncDjZVICrwe16G7ldvH6ljNtDTPHkUaxl6cunQ61Y/OMqYMjwES
88yRY3KNfMtk2+NZW3AHgfnHmAzksfZIhKI6DUKBgNk6VAZxK5JkZvbqlQQj7ebXb3Ylvq/RN6dQ
EAA6r0C3FlJNX7nZTFh24lqXo98WtNyDjGWXVzLqKiw6vooQV1MgEZBOpVIiyfDDdZStaW/s1tJn
b9LCEKWd+tMMW9atono6CA6/duNztAhaFjvmmNJKTDzYnqYsKc9KqLfs+aofm/hbiaqFvjz04B0N
B1NtK6FDq5YzO3B2BPD5pdu1zl0x3D6Dbo9L3DZJHAwoERcxiwES+KyQku5q2KcIVri9DwzDPzWr
QHO6IP1eO3X7OfDGeCMJ/thV7ff8UF612BcgHoLWZNte6veFGGCPPp0KUF9I54xXJsObTdTJWuzG
mVW4BTKs8/fveIRmI3vFuXxHLikb01TZ41/zN71rWqgGdBphZ4syPaEONS/SGyIMI9LaD5YClJvc
GrxJlpXSvlW0bi+I6m61L+IhXWcIQSvdRI8Oiy4CDwL759TABzXck/U3NZYyPrn2cYGI2JUKzQTE
Ejrgeu65uOK7BZpHY0vqzDfUcUVH6SooEgMAn/ttUl7jVG/QWPKXxV4fVhIBHZVqPN60MbjFvgD2
Aggil6SonqNcZwrlCGGb6g86e+e54RKNNCxpgTMpbRPxnyRQGwoI+5QgnnO2ctnfu3CfSdqvwWz1
MVNe7jYMi1Uz0uMCHZ61LyuSamGhE9C9T4PSysDv9z8F92LWl5vGxrY5SRLPxJYxtbeNUXAOoOoH
yBAotYsFMfFleaXlaCem7BYdr/91DfFbF6Ble42qnr/ibgpZwvz9IrKN8lNae+yERaiH9M0QKPaL
ap7ig7XGdwSHli/hliN2h/Jv4C/RQLCF4blq7ffUtFYr6iQvkvCYhW0Nza282uO9MVXHHFXyavIZ
WBTmZ8CGSXLwEpbOYZHIXPx7m3rU+gC0vHZuyu2EblblSH7APwxtMKzfA2mWyQfLCP0BDO62a3Hk
CutWoNemzOwHLKI0X4PVvH+FN1uPtOV2E5sxZVTobryM6nrmr5fueOWckK//jKpVm4YvcvTYHILN
m+OWwT/JTJR2j8xplH17LuSt/tbuZwbzHEe44UKO0ljrn/C0ubOyG3R8pKHtJSFGOkECD9Fv1kz/
U4x7TMzR5ELN9gx6xmLwxadXyctGv1iF3LE923G9vbjQqLpYWvx94jOfvilhvgHvW7alwboHboHr
csAIC8LV6aRftX1vysjr2JTv927XWi7ae4cpsg0Oqm8QGQuSw1ogjOSzDlv1FA8Q7NT7mSgpuQck
L1jqMuSxxuC+dJrGvD+gYvX02D28nxT24mjjvVxs+Gm3zbw/wCDAOIAxVUY8paTtAy7KYi61Twap
qYBYTy5zBY7i+WklITQngJN5AAMalDhBN9cEQb4tQjg4ic4wX4UeLVW6QsmyJwy8PwLfbrni8hpb
B+WX7i+Sh/92+KfW5zj1V7CLvxu3ZTRXrcPqzb9vxVw4TzlDrMGytiJxl/kM1+5OTU4V8R/WNyGS
4NzNEzlgBjOMH/+rvWPidtBqDKMdDcVNQWfpdA8aUk2NzFRNPwcfww4LWBbJAGm8i11P+q+nStBd
A2tn0Bi9U7Rf1Xne6Asbg+UP6mCBrHX4QZVqS70Nlos0ty8bpIfuhJxTem62oMAJostkPzrcCoS5
Y+9Xe+uNYwYxTMSwAhWI12mESSMmdgApj6aOLRrOl1QAYLMk/Zombqcb9UXpcYHJU23odcnjmRjc
cserD71sRwiz4fhDRKXeU6223PCLIFdOXdtDczPGgKC6OCmXOeuc/jTFKCr7UDV2tVnL5XIB5VPf
v7FYK08M5sKo0BuU116L9lG10cDU84oYo5j2ZUnm9uFBJBY8kj8dQbihamqafSBkAvV9zVDxsI+L
558y9yQV35biYDMEr/yARBJMEgw+hb0/04+pYm9t8LdgmWy/kmItElNfQqXF/2XumDQLM2q2vPMV
HKGMb+hLWoxC5NAkPyYnzvqNtFiJN5dofZn8HX7ql17pMNEQSUuAxAMq4nOPuPwiHiC2jSOPtBKK
xhHOb60hrUgebXAM4BrQZtfh3/owiS9ahVD4/Tttb5gkXVJPMXk+dURrP3rN5suOL8j59zDHCkFA
MEirR+IAP6DA7u1JOb9NwRsZXKkDu1gDJNJrLd/PST3R8poJFdGHVoxQYF+FsSdHIhgKVsjCuqn9
3Sak87juN+WnU88jqRER5jV7qoxIaae+I1ivG0DJ1Ug32PYl79gT/xvVCQVQomWwr4yhpxnTX8Oe
WXLuwRX/W1XI3bV1UKUM0AVLB0/07di/SH4qRNT6HPFU731g3Sp4idLUIhnvjsARFOrrPcfTF1Gb
8QAP+0gaNhDgaZyatPLAxh1WgsYLRBgG65/dMC1+Fn63JmCuRdfBX+WcyzcHjz6uasqltCX7A2kY
4871ziKR4q3y0QV29sW/04+4csNHYcm+yfULpwG04e/fQatKNk6aO72G+8+jz6zPhIXvY8Qi2e/u
3+S88F3bcqVOJNGijqp186IibrHfFdvTITVK4oCqSMf2MnVzKzD7oxczeQKW7562CaJ016Ju1RwE
yew4tpEkulSJMRVbuSnb40r50Lr0qaWDTZfFR+rA81PgXuggWMYw5IZrjQg++qqupuYAd3bO6lB5
iLc9VshfaVTECENS3i9lyhorPASi6fz7oSQd/R5kYFbntl8hW9snWqaz+78FZhfrNVffaLDFVDIP
vQ9KWOtDSLU+Xj3xq2Te84b/eqYylPXgydyEA38XGVz61pEzJ+mDAajhJ7HumzPFzOeO25GS2pJX
VQmN1fqG5Mx+M3AiPE7bUyazSzqERJBA0ntIIakAqfOJoJrMHNp07pXQv1SwwQR4bYDP0OAfFiPq
yOabsuq9zRTwBn98RaGZOVmRycwWx/hJitrxN5zZ2XJa8f6+7lXxNwxBmLLHAfePKTTdWPYhFCOs
OxZeXCZ34nlMoyKHIfb2VM5cq/Y5j8+/DegNdl4jv0ZC3GALZpcrOH94rqdiDR7NFYbtQ9jU5gpV
LzJiiFSWw+3stPhjzsY9dmkFhwXSYAamjBx25kdV0EAHDLsNkGIOUEK+/Pv+gNRZFfWHqyHoAqzw
PwD7hzJfhpJGxOW5U/7jFoJRB5ee5PlPDr1fwKL2wSBaCDJsN8We5+pgM2vz7jr8LAeE6AhJGMmx
b2xH/iNTVZ9FZC8hzb/TT+F0CwCAgh3QnusqZoOkyvvD1dxO7cwZ/BQuHsVRpR+c39LdX9KuQ+Pr
hUgUqTltVoWBOwRD8YFs4wb8bcnF/2I0i7X++hBTzQvpttJ0hx2XGkSgR9cPqC3d3YeaFhkhG0Z5
dpFf2gGmO6SQK1xE+FuxFVkm81vIGOI52+0FeJtmYD7PXcLAwSrBKsRbg3ZqOdS15KCK5pSNTkrl
LvlFCcaK7dJIgCrEPb/13uCpGIjVB3w9TLdOuf3Sq7tVQR629y9BFH+nfsRatMiBfP/GZZ8kvLxg
XNHEyjX4ujlvU7USWlAhjU2OzxdF5QjAwwkZRUPAwX0J/jOfMmezSgpmP+3retnM/DkZcx+CU6ol
OmkvADwSFiQM6drOmPOWyrzWpK8Xp/osf+HdhKQ74VuSiNGPUAwwi8FAYF8JbYeMIhBSUQZDkExY
IkAn93qbtOzH5dBCDHknFXYgrgOTs9uu9I45xD9E//pQBlJjN9FI0MhYCAhgjU5UbJBdLD85cnlk
lmVbQQxLPQvvK3eXhMQJWc+Bao9wFKTXxUskOJoP4BdztscdBz0UsTRKX35Ncgcmtxu/LKSu3JvC
WlPk+uCJjUIBLCDVRTU86RbolFLFJnCEeCB5lHLG0IHOkWlNvUqhAjOzLutSRu1zGRq8Zw4amHn/
avWf5ClGA8wwSWzhuUJGQoWUY9GkduIUAVJVjNYggQZHQVg22fhIkJHPGHnfGnLPsCAc71UL8IjR
7pQG6U5ljaO1Hg6fPcCOSGIubw1zyEhAdDKGRMAQLsRN1VAKb7AJjRBY8yEOnrHvTmlCCFgyXEVw
wUKxdVRyL6uq5AmVZQjYVEh3T2NUDmVuUYrrQwyzcBxaVjCXghJoMB++CK28ILNvhUIp/0vp2hVa
oDsFUd37AyX2Mm3wicQDbnu08CUueseRn6iSyvjkrsyqIfKP8egK0NpJL1nZiIh+GWdH4LqPrWUU
kYIhQ0vdiAip2hEvD0SGVAmAIBvs6DUoMZS0ySbE7IqQuAttnwh+afAz9uaz9a8kDVtwODuo7EEr
zPTJs2h+MvBFrbmA2OCNavEPu5Ymbi2iBsw4Xweda35uuBvVDCwy/xK6UbQhv5esF+/Mnef6PqZ/
2C/wPKzH85zhjJ+rnWgpGFupPcz+5L/WfW8achjRZF+6PTizcyrfHur12TDaZYJ36ArGMbcfE2Il
fCJDAZBbvsQ1ydEvtzaZI0nL9u4ZrtdfxH6OYjgVT7n1+P/kUWEddfQ8/dg5S8bE9wbjFaAjCy3Y
SqNJTVTK6k9yINeB7zp3VzOt7H1V8hQRYaBtyqwNv6QxXai0KO5PsNnIg76Xbfu5HrrMRTc1E8wP
sv/gClkROL3Q2liaysaLPdjJ+hQkKtTfe5bemRs4Tofa+fVyrjpdH2YSgvAx1VinlI3uxoGRZLIt
oxbxdQOh1Ug+WNnqE7b+wxSgUcbBgxqencD9vV6gvVNM1jm6lbmgrcazxspFmSBQbGMOCwNzmNmJ
Twk3nq5gR5lJy9yFc94D7ZHkrGnS0oaHLBQv6BWCKBsoec8hHPiLQndcmPQ5lJpS8bpoKu1A0yIZ
a7rXcuw5518idOTb4ZChLZhQeDnWqdL5HPP9EWNQo8iJFvNnLWEzyPor0S1J67WTkP5fFVasrkF1
3qkhbQwXj/hpj/uf0I3dBFJVTAzZVpqTN3BY3ptUtP8NvI8B2VZiCDxDcD1BEOXnzODQVo8fek0x
7L8Wygv8h3TPzX55i3UfdcIbsgOyKK5ZVJIsNrANMekWD5USvY7wLwqAFnu7smVa071E3ibTZ24h
i+Az3TX8Fd3SX8uaEw4qSHpRjAzJXsu1yhVOCsjg+oJHyENxDfgdrlPZW39FPv6MKkyIovpN8Cq8
+VQrE41+LkHwpSn3IgfMRbFIqkVYukdK0bWUOuUfG3L9aQTuc/kvCrD0VSc1uKVuKbfQwvTAM4mY
06rdz/e4O0yNSzL/9Nd25imToxa4QKw4Sw/yP5m4oouCKzGuei6fg+B11//0in/5NSchkVk/7fga
maIZHjjmEoHuJUUTjdhmCTVMOcSberx9OJJWYeBjkdATXpB+RDFiboe7RIVXKL2Nyobz03nA/Fnf
Prvhbx52H3BE78PTAiDC6wbSlh9FsoXoDfvQCcOE5sMqrhHrJYrwMToysowZs0YdGB8aFVmZXutW
92RgbtddRF6KXuDh8bMcBEOAg1yUV2t0kP9CCBviGqTwWNoxr4mjrAhBq2TsuGqc/wAxgOYj108P
Y7Op1xT5SXZh/4c9llSmu9UI0VM1FmZY6isMyVmpwwR/8RGk9zp/vd6lNnxdXOTYVBqJZuzASRGt
4mVGYLJlKNC6ASEMmj81q2CjmZ8gJXvP5eyjoLpMxUdg1r3kyg7gJ6CZRtAUQXa1SHkeNsfpPrP5
cY3Q5HYLswkbrgN5ZMrI6uchFlRavW9RLCpgb9kQ1tSWvDPJj2kdtmUfE7tnSeinkp+zBJQROJax
2IBmaHc1+2cLmHDEaWphl2wVbzXp05XWRTg1S74xzkvjPvIDWYzMr0Y5OkefFULteMWC8uXrXkCo
zr2Vh3OGvAFAfcln7KVyhAw10xdE1QgSXP+fOxcHDQy84HNfYsq+YCPJ1wj9Je5ypJKJUdX+gGYL
k1QeWs1WPsdSzkOuJlRm8vkeMvxzNXxNaHxUUE85nxR70+PWTzAIPNRSozbHz19EddFA9CXco6ME
oPXJEKQ3DTDi4Lpkf7MKjPIqiZ6kN0j9uvLblDomPGsEO3lHp+HkOHez+KKzoM0BtBrSGeFvajnm
M2wH83wc0HvXbD9dWx7PuQVbplBaxohrzjzJO27l1ur/PAA6lH9ju7AUprQ3l+Ow4mBekvq4u0xD
Wt8nR++AnUcaN1OHKbf4FXBPGoMPaXhTukJsxWnlo+OgoWkMC++YVWZa2FuMMonTvaXGnlK3OJdY
n2q2uwggHKqY2DAgpoVYHWU6TPaYWW0M6mxwNGhPqI3UaB8L6tTkdRsLkbQ+P/FXzUeEkIhWGr05
S88trZ3iZTlPG1i10Peridd9ziVMRYtqm36pdORD/j/QCQ3TTWZLpDC9XBdWsW2NWVNSMaXGu2B2
UxBpVFNO9pCaiyb1ZjQ/jD29KUYoXonuaiaD/P5JySlsZySW/y7d6GrXwdtGiZamp78ljm0nWD/o
9qUCwSOnVE+bjAB1UzD6bQTbqLuRByZB6E+TYCG7/hZ+4buSk8KzpqY40Wtrs5g7zOrusjCZMNUf
jqQ2E3Vl6zaAPmBTzT9dQyGBKsuu0Xq2yoB/H26wIemv2pejaYaUH8f87bQoinJ6q45L8CHvjL/2
L9i+NjR3eMgwBIpt4+xU3j0A0e2+Z1OmDby6t0Es5OZyqj2jBzpeXAPT617RXIoY8nPEPgqrsz+f
pi0J0qkyvkV5DIx1Qt3yZOYlwwIfl3Gngiwo4geNWplw2HSjpJUU+iIV5OG11ys3iMphPXrkm+6c
pZAcUFCpZYrd4q4hEwsFMMIUc+Lrl6EEkCjafWDo735IFRww7TXiA6Y37GT8xk2cjnc91Cs6BqGb
bjPGzjPg4PHnTpKYGBEfon76R7q7XbTfGbIeAKhdiw2V1CC+gvcjZPlyeMd5Eo1CxzlSwyBm8lWs
hO+CiR1kgLK4UMvqmZkVV/vN6Taa7kR+E9i9ihe4JouofZ/Gl5v75HbpxteLsIZiUBB2OrocKRBK
4Y0A+K8jf4/ZKbQPxkjgwhpJnc3MN76a094SWl3DrgoacP0xP4dBLjLpacsCnklZcBdqsBjsi4MZ
TwvUgfmsRz2qnyMUFp220e/pajZEmjXzl4q061Vnu2Y5M19xM0VBi7bXtG/zdks4Cbt++al8shhG
K2tEOYhrUwzCJe2SHxOSaTR+/xdiMNzur3QHpHkh8HfenlGf/UoaNb7+Ut6LGbJkQNLekjjoQPUS
8IvRDdFRdR1CGsgy7tmG1xCuNvQYrw8vCVOowQifyYiJr/TBHDZs4uUPlZHF5D+njh9dvpGIvz0Q
sex/hQuR0M4pksMwbW2P1L5JtOUphWN58r0EGr3GrbYvd6dPBXga706iNQ2vqJMTMiGJhqMBrjyL
rU4q+AJ48nhlHT8JvGFGySDKf0t//iFjuu/+nBlc9QGc0kzv8aClTSe4HdMQUNKhBKJTv/EEhAtC
iQ63PzrJjqBUqToCA02igmjLz5y0Ytg+jcbai2vRFGi+V74uOZTv1kFlQEXidtZm+S6E0Ym0jYvN
S21HGMPRrQ8Iv7mQ4qZkH/I79gGYBOngYvuOD3EhuwilOY9copr2hUg36jV1aw0k2/ACFmyRYMrR
c1XopGYN9Dn/Zm9O6RY3rsVyxpapIvHQflRyLKZF93HOpPsHraXxnvaiYgJR47sQ/8GxEJUsUB2s
rpDsG129HKtMXSIF0jgGohk3Bpz2v+4rVEvVDjWY+bnPJsny5lRawcCAZ+i5DZyp/0raQs3HxfAd
McPbk7oVOmDjEKLRZcrzApN902XI/13HdEEIHfg+wp10CGN2jCGT41tFce6lHGC0i+sViFJ8FsBc
+1+Kf3VjiGnhKK0l0mmw71eIBE7RhVahhgY3zl3vBgU8pQmZAFm0WKo7FDkiFIDcT+wI1fZqof7m
Cp1hd4AhCK+2uLGYNq8b0FjtiEbdWgxwMhQsJofyfkcpuriTUcG99K+sr03+2Yj6sC0ZSaTjLp5z
/4JANHP1MzhE8+pkDUrtQVvBpMVXPqCLIfkcZIZOKtx46HC/flmkYQHvVhEVGCMQguoWCvVGFfrp
6omN8+Nry37ronymOJM6GTvtp17NpL8Ly7lVRSlFqthqO93TPx9Voob383oYhCeg7Nmjzc2utKyA
QUqoeoRZrxn292JuAe4bmpTmcnaMiAka/QI7WYFrEYNhsIbOvNLYfkpYYiZnK7I0Ab//ljdMvwrC
QsQoho/75ttX0VSAjYLrHLC24d4iWDKnNr5a2WiQ5fbn4TPe9KQHUnbTfaq3PQoOW6EC1hRtmXd8
NiHN4D+KXDbh4SCHcGWzIkIP+fhxlrX6NboCvp2oQeXmAX2nVRaKQGeVyhVpqyZYM0KXuitJ6+4C
CnEaNqiPL2X2cU5wMz2Zmlw2CxWtZsVfuyj1iNc5HjOHsaDP2SWfiIIqY4IZ22h5VKP7aCRVbkUq
Yk/6ppOi1DxU5nnR/OWGXkU/QRq09xJvYpAlFWj939UBveol+BNeRO/8NkSOmwOIBjcb90MzDaGj
5apgXv6BybswA9zLvEPiqktXT3xsqjBN1Yt4f7ht0+HczX+liMTaohNhFVDSGEImLvVPzM4gOi57
x6jFWTwgUganITTV+ifm3BOKxXPXk1ZMxZMaRQ+L+GYWw0wYWRZ6ZP+pUQcKkejKWpNGiNHxEGaI
qwN7tXd3who1CP7/FKDceJ0FVJzxLmzBC6Zfpd0jGyaWKtI4+xB5HWVBrYivAgA2aBpuZqPZRHVn
a9MG73SMp3qtpxz3vd1kB7CSQdYWkNL988xJWmj53VW2CXyWOQPaS7fIhCNNheiX4wSZZxxWB5fs
RgHC1342x03tS8Jqjny+wEsQviZQaBtYcCL70qQGCtnHpJ54B2jd1q3aXpnMvGaS5Hoba4dYQM8o
GdVVw2LmqYlechpP5Hk3wfBskBCmOMnTQEy//aPevO3SKrCrKntLJoF4OUyrBRsI6pHeKUH+hhg4
UbWrymWp2BpXHsIs1pKWT3PVEvlSNC0dqrnHYXC2Uc/cX1vCk0zXZdGc4beRWfqeLYpb+sgKo8AQ
e+JpybpMNEifX1u47xwR3Z60FAxiJBJSWTYRP/0n1hsYpmSMaGfYbadt6jNYWWEk5kS66oD5PTAX
QysBG+QZwquxBg1Eb6FU5ubMQWGzBZFRE/4aN2OPN1fYu0wlrsqiNvPEtULWjJbORCdm5uKtRucK
DzaFstTbmyH7V81pW4cEHmGwZIbnr6636F1INuldF0w3sfCZQ5HIkFiwsFSK3dqtEAZtrcfznZWE
0aUim5GyvjXT7Dt/njZbsBk1wz9htN8dGUHPa9+ZKBjitJtdTUfiB1rQGIe2k8m2PZYHbvfVzcEW
oPrR0gV34eSEINEBQVRmu5AtJOSEWEpcUhsbuCYJw1WL2Iwcm/+udaTCxps4x8YooEahMJoAwDLu
UFrHgGtvY2cFbCNTw10h9Q9ku8PUd8Nrx56mgktfps9MeqCPtCmR9VYOFCrvLTMQc1SyhOVAtE/l
wiV1QWvVPYCXTjKN7Z/y6p7MFPH5Fhr48uHfMVpja2MJvIXlcQDmCHsl3SqoBYmU2feeSfPlXhh1
hbC/iD1hf9PFVw4Snz5h4TdfPsk7w9b2HdDoKv+VIKY62ufvzPxGQXANtJMjKnBO1Q6xoZpexCGj
wnQACUw94RwqndEmdiqsoMnsWMTkU9CK4wpnSntYQFuDAKimmUcQpqWWp46DedQQYV1s0IpEbkFT
ishpnEP8DqjrF/a4BA3kQrnmXuy/fKigC8T9xUOUf+K73706nBtXgsN7XJPQn/QdUMx0nMMp8d08
oM0YcQTbupj9Avd1ppe/VgMg93BCZFBTEheppBosS934tlRZ6wx9aacBqkzy5Jt8BPOyrrADhAcm
fRk6B9H1tIaXyCG6Sqv+klthKPsxSqB6j3g7QB75X6h1Z4dCdHLfSJSPBKHpd7Y1Ytw4XTaoEYdg
fvb16TEDVLGJsPFK26rdaCsS44qc23V1Hl6YKprZoUso0S6Nf4v/HFKIt7EbiqFiTiNAWn+83YCA
vGAknTydFMSkDM2dh3IMlzN85NEaHD5V9yF0xvYaUrH85NMV8IjKX7JukbT+0L8+s8ANsUSbclIg
G3a78w2Bq91iz2TF8pqw6zX+VPOVWLwr77EMf51jEJupIieBsC9GVuoL9pIuXR0KdSMfKQf/Z89D
aIFMKNJ4Z3dySmUyrPi56cWjUwPqciSvnMv9Hy1D4jbt/7Sw/dJVcjlTX5cZvX9CDPXtOcR2+WQ7
3QnUOTObCJTExj8OBL725OkRDYA+VSkQT1gGMiUyuqglwndrbDkCRmChyXsoozUb4WJJ5LBlLoeb
ZHr0Reh4zBqozH09wjK6IUZPeGjblle902fYAxORLmNTYqzQhht/jCwFBl+T1Pv+ca69Wbc4onLJ
SKXz1qS32Iqo31nELop6O1Ixx973j106/aBOBS1eBDKZmmgCNUkmhSoD9YRmKG13osTiXoj92igK
4eeMhS99Qr4Jp9gwV1CzVQ2xXYcL74rtbXrKPcSi7ofqGTnVDvrErF+nBPQjkev1t95ldVurpTGW
wjsHtzqh1sE0StHsqiTsDxnNmT+IBFANqMmJwi9m+ImJTrF+7wazEmSs+aHmOi8LnqXRGh1h9qcI
zQ0LYcTU1quoBGBJjXbWFDAf0XVGZiADHhgxs8yQ4hvQ4RE2RrvXFbjU0ovk9pPcPy2D2jr5aThG
wu8u5YjL6e3lynqDX+oGQ3GEpxK++JEAkPAv6Ik6rntEXS4Un3mS4tB1pNCIbnqbRz4H050RklNh
NbC3j4Qt7tuzLNa2JKmP2+yiX2diszfqcJVmzRU27ir9wC/4d8FNKtfRETwgPcOroNzQfxZWi+Ca
gfpzBSclUN8YZu6LDCCqC7/TVi9fgMZsbZ1Z9eYousdhCjYD9b2sfmnoLB5bXNB2ZfdxxzvMIjDZ
Jyobg2aYLQUqKpeLmPm7xhJR/u77Q1kOdnBg/Ryra1KKn37ZmgkeXQz1ZROpfdyF6DB+NjM+K5Ea
FBR0MSMEc4gAiA+yYIoLqBaQt4W+MT5GC8R7o5QWX7gyPisEsAwZd75TcjfIgZGt8WI8ccUDqtu2
4O8WAk4yZUbVC9F8EX94CNu9BzIOu8qStFyCqVpJ7jVnLjaoW3K9dEGe6p3ztTEM35QOjjXmY/nE
5rZHyg3++LaFDjwt3rXTOMzHrh15S8N9WPMdSveU9/+myY79af7UbKXZ0LILNUqmggVk/04dLjdc
cNnSdDtLmkfpjPVZ+NLbNPrn0NQqF/9vtlPx9s68hjKXXhKGtFdifR8rUXnRKE5NH3NVdEYH4TiQ
YH4Pv4bLZEVgvDG9BIFD+12Z7brpplg/NbCDx42bGW8vwJi2MTTC8JHeZZwXA6ywyfySsJR8V2GC
XqVPXkXxs78hudbqKFxjzhwa3l32p3lI027FmT2+Q11/H7sYXcnlyUWfKv4kBmxp0H+tloiosUmM
ajWwSZd3oTEwI56U1hMSnh+irSRqRLdj/IjF7IvUM2T9+ERtZOnLGPkx+xvj0G9AvK7kNtNy0JYH
KYutdEyNH4prAxN1PxZL30sNJgbfF/K0Fn/c2j/CC+8IeN8R4+3tbgQfTOMaxOddk0ISwVeZj3X0
WCFGlG+jcjumQS5QaAZe4UNQRXfm+OLXxjKzACBSLHB5Fq8DDSJePTuJlG2oDof5OnCFW8gYOwYZ
KlCJ/etKwhKTNJcvzpNeVdnPCGHdI4JDkIjAS1NIP7JJ5Pg28S8jsvTW82J335mcnkay50ar/wkb
EYoWr9Wj1tzxDNallSxK04UbGGnEw650wcTRWkNyxO4EB69b79K/Vu+K1mxup46ZIf+fnVH/MVZz
fr5S5BFmeWjwYwVYnBCbh8dU2Q+87SsPvwe0+4QT9IHcpqAI9P1JXLKaZKdDqrxbs/ZDOJpEC74x
iMVK8pzeP0bLVOAMINvWoaGaaBEK+jTGsY7AZZpcLSBPUYrqTaqGpFI4BoiZZ5/eWtG+bofQigGW
jN6+1dDAeo5yar+4bbKuKt6Ut2GPDBr+vd2Yzcz9azDrqtaQIawP0GegpxiuLGUWJPedlBg2bqxI
SFXm4qndHQDqNX0KvM2nKRjRXQ1n1fJRkx7D1QbVR3300Q/jLOusiN/VSKkfDK2vswqAfKUnZnh/
5LPscqQc+n7862pJz5XrNHmdIz7SaUSNTNIbImLJ9g7h1BIBVYhTQRqXarnGZZbRqLj+m+MLkI40
C6gx7Qp+2LTQYu6n1gdRQSugtQolQmaMDlvl6GiEH5CQTbakup8tV2pUur7SGkfEByEGxEuGyHvX
LaP79Fly0ahja+MkDNmB8rnu/54cnOfpKtXfy0nvTcgy5rFRs7QjYd/QQGIfmLEbZHOUCm3rsAEQ
e+MAVPCPLNBGcc0rusxuG4Kuee2ZtRDDjSuubsO3HMoIVfUKylAnHyLj+kTwY2qEoSu3EjzpTpd5
W7UbPlR3+MX5i963WrYXUm3razf2qor8rP8kBO88pIfEc+DADIzX8WIxEOGnaIw3C9LOn7r+VRNX
Bo1NNHtAht6is6huH7x5nDIKsFBJEd3esPz3Y6BrVzuOh3//VUFs7xak5a+VcrxvP4T096WvM5/i
llIgAILsgyquNmXi00/tIqYGrXZFz2ds8pjg1xOXv+xouCSrq4Tj/kT3GJ5MIJjn4hrTQZX1zHBS
RKIZL72FuAd5IOwem2glA+jBUfeVPtwp9vv+6p89WgSl8kqdek6ziITXratm+N4rrdbwqY4M3DWJ
EaIf8Zsc5TlB1DhNdiR/l2rtAg4wBDSDAQCtrwV8xNHhDFUwTwXgWQHLAfnyI1YJJ76uAuu0jrXv
svj0RSGOcEYQRiPozTP4hclu06q21WIhovFdQaFQHtpwsLD1r0BWvR0pyrGBzFkS7jVFfxSk2m5D
38sDKrNeDh9O/2KJX3yDHfU95GraQeOvET1sKilcJCIxwvst0kHEp3oaZQih8umHynsgwzZvSgp8
l4eOZO779U75lBetSbwH6XWVd4N6fBFBpU/jJ4OyrE7sYsYiKAxiKgFusBCTAopW4Z+aT1BPSCXj
AWZBK2ebaCj5wqEx2syug/HeuZ5DQInG4i0tN6r0DSplgyCiBWsV7tZCGr83Trd1Eh/BZHUVQzrN
sbSPy5v47thb1wS8X1foKPiWf7bezUkWfc1RA9LUdcgcybNbQ3tKrD5UQwrkmXzjG07uXshsixZQ
h7KXvmp65rQ2zALFBi5jIuXO01Wwh6oVJUUatbWasjA35cAzSL5hOlGjISigf48VznW9mF2II4kC
5lSyhBXcSvpjWwGd/6Holid8NkA7gGJiLP4lAHeYrRTAkYKpBsV2nvb9I4coRB/ZeJAiXapE+9Il
WV1pUuTYUTA+En54DWq+Ei7rPAxC4xe31kLl5Iw/M9Y/ai9Cifxc7aeL3rvnnk6XNCsttgh62DK/
RRY1/UuKypSvFHdEAtGK6wHl7zSpOXtZqoKPzqEcGtgNVErVkugQjc2RDdY/ubkbYIow3j1Q0wPm
Ech5WshQ3AOzF6a8a6W1m0fNTDKG6aif+I+BtarEHzqrpUqO++uT/liSV9fdtGyGCHneta1ou9/W
QffKSRXLS/X+Um1KqEVNyafMg+EnN86ZXhUF2vE6mGmWXu5i/7o5rAOxjk6oZHfjAInItAZcX+rz
EIis2hCBoX8EpfXdno9rG1+yVji0oDJrRLjyphruXp2OB1ZdrgMVVkpd7VtJMmwQE5NoMcJGgI0G
msoJamx1AgSBuKXKi8GndX+dHEoaj6LOlxuYyTSf0RbW/q0PmtDrzcjJAnDV1HBWlI/2ZUEPDvjR
sQgtTrAp0dMIS7AVr541gM0NS1TSm3fDg+utICOvH9WmgvDBxC9EXI/P4KViw7R+b9iHqS9lwUsI
wlkC4XqfVpnsmuqRleSiJTLC0Do1gKNiy4NgQ+g9vg1vcwSWxMho/L6UQV4TSuwfHaM/GbVaAlkc
49AwH7/lvzOBTbgmCaURbN1KXL0KT7A1q8U5oq/qjn/2tfTCYaXpaTyrlQUDMfDj2K5E7nFAra8D
uolVz4lGGTm9qg7XC0spg/ZH9p2mcjJF0ysJN+oXjUpoLXYTlYlKiVae3GGM68zqfkQXfOQlOsId
/X1niFmtfLIkAatDJfgNzfQYUYorKfK6L8Msjnu2zJEGbpG+Q5PkcyG6Giy6xR7sadji+K3YUFT3
VltgwXr0zPPLplKfpfgW0Po+Dgh5N6W2bwXPENeee8RNr9WeINm79e0BXWbkBSfIb1IqetHfQijQ
EDi1aSuw2KRp8cQkSgmp+Dwq4rge2bYlLSzNNymEaBMI4m5SRXpl5PonbtGq7xVppZ0c4s9amasO
P8WufFLA5727ibOY+gSP/s0bASYdbF70ScdH4Taz23B4OzU8EE+65VVpfRSycHhwTqMhDw28FMyC
EJN+x3fKPrpmBW4lW8kcho6suaymlK8UQspZBaBQ+CRyq+7B/sDQsn9CMKOUbYd/ciRDwBCZSPg8
JvZMdEmbKeve5U08F2yYDLBLBEvj3unNZJS4ZTjcZNTpkkuLmjpUzQva2ZJvvF+1Cdz6YgLEICt+
OqIs4RHtVeP/tHJGclQtm/wc2il89U0n0MfPtnkOUP4eVPv7Hxm0+jM86RLzyknNe8V1ZOd/l/Cs
sVXht/9dUTwTllr7oUb5UJ+WYksU8QFHLHbJGFfWkwSimiDFBdx/6fCKBnZJq/IBWL90b9c017oA
Uodx+abnx1IclKHXq3a006/uniGJmz9DyyfbWyfWHg4EyE4oHq1x8t0ps5qqqoxOLb3LhLjdiNgw
BnwZmxwqsBzioFzLlGxA4jlFgtXybxHgJvAcltNsZQ+pcGPEkTSJThTHAKRfJy+QDMS4/ATyDOpF
KHvPVw3qze3ifuz1SWH1Cl7YDxcjI80c0dA88hZdTptGbWVUwJ5b0d+HHprXbREFZwuQ8+eMSY6w
NsmvVkYFjJRA2ncu7pK6CqwlY38l/UB6Zb7+NlaqWa2UTX3FaUAad/jaofue3fLAfBC2RIC7+V81
jx02mnw5/iFFHNCeQyu+BkfHOz2ORu1frC0wUsXLF6hrgcQGF/vFsKuYvabNqsBKWzMKJzPLIiM4
17swHGY3P3CHoW3kVVaega/cAR9+daRtr6m46TOIuRIXbPzSQEYgapMTHcbDOWqQp9kUEis8e8IB
7A7yIhEcCQ7LJFWTREorA/7FOCv1jJv+CB6SboH0RiAe0JAR0JDKQZ6Lj8hFtFJ53dkuLJWupz10
Lve2POSApp0Vw0qYn27ELkHjonxcMdeyPB8JjEiRHiOHFD6+6b5fYInpCi1oGrhzTtdTKxdJerjK
zBYaQfVBUvHRY2JZ7vnvCFqwn7gnqpFN27hFtFDEqvfHvh7mlk8TUHMO1FxuNr4kwTi+QdX9XDd1
90isIklJUsfaco5DYgPwqnEbhwBTd/ZBJKgJHeMVRsLBtMGoT6Myp9CODmRJxfPZ3eE754Ibh/3b
psSF+n5g4YgSZDFFPRdKSQC+QBDbuDxgpzBcQXCjpA/SdCEB76OBlGI0DOUo450b01vP1elGQdcM
nnSDfqQYfXgUeSw02WHfPbHua/6lEEV66FRczHuIrXUVoFW57ezVgRhUB436vlEz59yjk1m0b9JO
NpDKJF7YxjRoFN1DLo6FazmuFJtZRijAqzMI8sqOphWmjF4Ylf/Iiz8Urw8yLLXg5nMIyCOy/xhZ
I1hDHPPlvnI/kpZ4apG5CaXIGTihyFH39uknjItDb81K7Yz74/MiNzYDY1ZcPXu3UwLisf9YunAv
kMzJZJnJ85yjipo5ovbYOdI37jtxO1O7j8JzmFqUJ7myEuujxZX/7vMMoSfDXd+v1mqIv+HBEAJj
tJ4qhG3je95YJ/OaKuZjTYWMAeisJLAGrBKku7OIOzHnVbE87UoyD1w3FHilQ1Qz7pOebTn0YxDU
LL+WSVcoVzUQcSUmWLp7/KB4L3qkOC33M0cKHyUQHL8W7cXG/zCZUdtTR+5R8WuZ759dToDUr3b3
DKMwRmP/5dovD0exDiia+lWBUhVdPM83R2wkpT1g9mZ/ghIogrJHD0+NZRmLw4Z/SDgDhxs2kAE4
dvz7wuCycovDW/bk+KY3CbKA+Vs2SGR7H9JL/rvsXH9ds9YEJlUljvylHRNWK+xvyAX2W4+6diSE
FdCx1w3qBEc+EDbyD7/0CSQcgt1LxlI6YNsvPytSy9lRYYo+i/BF6FPlsh1IJjiH3wtp/eleLBoh
1Ixznc9Wi2m57Cy6qjCefLtkohew1X04G6zfmqrzPl00f/ScstyNvrZ2JNBbB2Jgz1gvgfhEPrqS
c3M5t/L0njpAFnakLIqYZyOMb9oiXuc7eoWbr7d5FzSewQZWQjex6gTbOzCjDHKK8IcJ0Ofo8ZB8
dp0q2JyAwXLYPArk8qpqvwMvav6q/2kI2hEYBbKvKK1EeNZe3IXwNhc8GT+JIRnQqZMXKGgRdy1n
pu8x7yp0M5vHZvhB6udbyXw7mhtSG2a+SIONnqmCQTuUPtPoTTz76PvfIeKRxAAWoYPEEzw25hV9
sbi+PN4cxjC3v0O95XEQuj4LFdRiHwee4t4ZwOE/QDPSsTeC/Dx2AjnqBN3YcyZN82S41ghtQgCm
J+x1jIDe8rkrbrz8waYEPhNR2UCBtMeZn5ElHvCvoGM/4VJFAp+7fj0nKpeMuQ+RoH8KRsTdxNN6
40P3Ih+mEP+goCuYsJEcWEOJvCoAigGaJoGbhkDdlfWlyNT0P9fJzkc2Pxglo92ZjeMuP2deK/uM
ZdEJMgZeiCcHR9QHjpxZck8yhHCcSmh/dZTaFwQgKMjMxIPEVzdtSFQhJgC4T8wWoluvmqsZ+u7Y
AQQ7XQ4I3Ji/GonTBx0kQeziCSwXVjxOhyczir0xxHDWT3wxMdSdFFIiFKrNSUGLPImRZPbrsWZG
wEIExnGa3a17gBtsTJQEktqKFVPcogeKTkLQ99AtayWQea01+/FmpLqouFTC5jtZkT2wA6mS2ZH+
rKWu8ZM1JBBn4K4I4oFauvdkbSQe54Ned8MdXiBSWmB2DZne/cDsoQ/R19sIpjKoO+2LRv9tHOpg
8Byv38WpjRosnHbEMKvj8JY9rAELkK6uCBdMddy8qv1kf3mQ74V5itubVF0apqD/cDzDGnd60DMU
pi/GUmn0vDy9BU0xRTnGCpTOiiJuZ7Cc9hBRkrWFf0Kzw1IKGR2uFZkhUtJrSy76cKTtaaDSUWhS
bleBjoc+7iSAHDfUHp4ZL6wButNkPMEoHH8aT3P/H/4mPLYQ/hyDmveauYOaX/OSblkTdJUdNMcG
15Lsr2FOMB+2za8Fj9b0yfq3ewc3IyFiXQ8rQTAFyBVJN2OwRq40cJiwhM4ItxYdxu7pkKlVMJYj
3S2J8IijT3txk1d8AclAkf5CTSioqxDSnQ0B61TTcQNLS7VUagfpeY91L7dx0BY5rzwasiimcKVi
unlLWBOstpi2ckSoKnBBgXTbCLbPbwjvLGTSqZY5dAnZJOUMGyoYSGos6lmHpVuPHKCbXBE39Uh7
ZHhLQGzrXqY5N+bO3bToqr+jaZkilUkMJsEOBLc9yAprBE6zFdTSjzAW8xlvvg3OgQQYg4Sa9V9c
9SkjZHo5MEdnIQuXeNieIh6tZwY+AIaGgvRAMF1rHt7MuUE5tmtr5tV/2uWKD9Uq39YDy1AiP92a
Mj+ooF6GeSwZoDqxSHdegfSUvLRc6qmfDe7JpDNq/Wu1n1QmkeXwZy4Ur4llejMVwzzf5QUMUvrt
RDBV+R3KIftB+DoqT4oTK96QIY3pyA50KoaO5IYr83SF2J51Dk2kWV/tDXxi0HtJ++ttpxjt0iih
/i9Za2ZGOvJkzmW7X2uImgDvOTs0ZSo+XyLwiPNt+LBN/mokbLxfPh/HaLNGip4AeG6/7i05AHKf
/Ow51S4G9e2g0gy7cGMjUdCgtPA3j21Cd+zmvuSzHQPmlZ6t9/jE6ANmJBm05CwCIJRfn+YBNlzo
2aVoI1lxj29ALlzrFcTYTIZKP7pNolMCMGMVuucm+c3DU2PrKFPv+GYhfhWAwZD+UJ37mvUY1r8C
uwOqN6B9g5N1ccwuP9ijaTryZu9WiYptuvRQ72eGcdGm4JTYsaavshZXBJwFlWapLMoEIdG1LdeU
J2dBi36luDQtaZB1gnJc/IdZ23g9DMzOsQ++FHL4BfTFK9FqWN6CijcSE9ZSsHaeDssgNgt1ASPM
CRpuT/UoCeOtZEx6rZrofBaN7blANbyIuR9OnALr4KQmNbf3l9sqT+UeTgRJx+SnnXIco53wIUpO
4grxt6MBzzSIGOB4wvjHKjGxuCISVTdmF5MSDh+4g+OaKJHrSRdUErxN+Iz8i0pCYTTgql6RvuwZ
/Xi79X8wFi2P4vIkrFLtFM+qqs9ckivu/eqllqHc9t//xYDCG5THD1j+87m++QgtpOunoAYABvny
vhm+WEqn+ztfpn3hYufp9n2eUVK+Kd40d0Hqr64UgRNPlmUyKIkPNMC5CvCOmVIsTz/D1J1w2kPo
9Kq6HIAqZ1qh8fSsndnIG7zVtUIZeNM+3g/qLv8yfaeQGvYEltuJBfg4ei959DFLNsuiGYkED7sl
d/r4UQft4b2iBso6wcN2ZeU//apNb3QrJQGoawkx7g8mH7ZnCtFDyrgS7+k8BXedbYVoiyxF1iPR
SXSdeyVPwy5H5lX+tKJK/J+FtfR5Ws8eaH4nmDIyRZfI2hNN+F0IJcpesmJfVx/8uf5Dpeyi0odu
dPgNKNaOLZUe0mnmeUiyP9f0oS4aVPHekUYsrD5Oczj2d7rvpgMzQlsF1bOql9PCJXe+gHkMwLJf
kvwcMNBZ4dmDKj/81Cqbxk7M7Dl1HGWZMNzLFEegqpQG0AXA2ZtcOL32w4AVMLTk3RiWysDYUd8i
jaaHPc0uKWocNpwdApWHBynzQHibGjm3bWkGoOjhu7lAOhhD1GknZmSXg2lIJs3zQDZLSfcHazFx
bQtP6aeQpuXiyr5HLp36SGxEBNsqUfD2BfYuNwZnsCqVCPZaRDoR/lpW4T+vbpcTHz29mWL5jH9q
ED/Ibi+IKCVUspRpzNS1jxwAtuYqegbw6Ru020p8AvpeM/FT0bsVnPmtcaoPDJV1IbhnMaW1tEtU
05oXJobhY26b9lPT3GFsIUA6WDzZzHfcn+U1wyFwAYGntRokiWaTpgbNXFlNgPHQwP+R4hBsI0Dd
rDFC5ALfZbqTAv8x5B6+kaLAiEVT4BwAo+FM+aPO71BjykCHmmWWnpcpMZh0dVb5/W2CZ89jD+HL
8Nv9V8KOfSR/1ynEU1HmwGBvwMsg9z99W78Bw9JzMT+kCZDDj2XWVQh14pxzmI2oxJM1eDiruOJ0
sES6P3+jgllywR+RK5X5lBp0DRczoX0EfvKL/u/4a6tpg2F0sJGy0CFoD41fzWBgrGV9Rs/byO60
SNeAO5JPRGOweAEA2X/hmbf/3sKnHPRK+60lO09Ijn4xM1lKPujWncE56B3WP61T++/1YBRdw82s
Xn7IQMfANJ9v1TSdK4X7AmOJqri3Gxwp4Z/MWnxWDmpj1+qowx1kW1266ocrYjK+dnR31jAaJLgt
+NQMPLCdBmx3uCjrJTaH7q2dV2fonhXdWBUbp9lj67AKY6oxYH4VrtJfEhlzuykTP1F8eiJxrEet
v/H+Gsmr4hiYAYgFpLf4joNKwa/e8K1ZMf8TPTirIEetbTNwekz2X6Zi+dVIX1/gGnmeJNyTf5g2
CXgsnmzLsB7Fj7nIQZBp6/CHSlJPTsn8VTbjtOUqQmtXKPYCFGE+9Cta7bTXVR9ZaM9iMQpqt+nE
hdoXCh7II2YKNH4iXC+pEGV1ZFjJ9o/eVXKDxvKVAuIDAAyzcC1BNcvK3vke+wZw8xfHf8QOAF52
T1J0kdZqF7oD1WjabwZSS+vWRMaI8F5fqE3URFrqA8x+V2c34wLheZY6iFk2GdCjqIXeoujSz9ma
i8iwQyUyapRKQwu2QXEn3sCQNE95bisOm5zicLZ01sK0KWNvAotVgKrLopKVJ0eEnSQWNBD6NJDx
5OaieSAnf68VYELvkJJ0Z4D1rrlc/TDSYpvC4IHLDLLd0gXf8PT4mSz4u0tY+nH0HbpP+4qxCR/Z
awCKvoBlrTp/lM55x2v6vt4qNKywkvmKQ6bV71mxW5xlQIzf0r1GMvdbRIyrZFrhg4+5w6Oh6GGH
ZgjIz+GlR/MPUsMo1gc9v4XJgNMKlEieRThnPfMIyDoahG5T1ypdAtZwoFw/batPT7NnmweurV5v
FY7EvnQfhsyeu2BZ3/38YHGyYKGIsVazqe7QiNZrkuIVw29P8/9vdAdMA38siq9vk++lVQUT1PUQ
DDhGBfODn10fqucLt+u1hZkE1ido+H3RyLW5AvmCzVjZ3/kWjDlV4V4oVFYJhdqjUjKd9xzinrxH
0tInm1g8GdMVhs561L0xcntOQOSKXU4Hd+0287ud3homAjLfRvpgX35Tp2HwHT1lB4jOWIcVwSvK
70qPkGockFZwvJw5i1MUxjtV71+E26/Fkac0w+aNQ3pBJnP3VqWqQHtxKpPPhsE1oSrToVoR/AX5
pkCWTNW2Ysgy5i2UU+lpRvM4GXTlKoIqwVSOAjTA5RkGGXDsq5fPjnfvLZPKKEHBit7yEkf2Whwl
HsLJq4yu9pxn/xwSPi8AihW8Algz6RuLVn7Mc7xsRg+lgvesfWRWYMTPVCIJaQ8wmNG0xB5zBWd2
NNq/8uZFvE7d6ogRTZkUqfFLVjYrz9f31tkawMQAq7iT98rb7F5CfqQueCJvVaBaOsf8sBd4yw8P
QNAfxweM/9RWKgxvrTxC2rG1AyyAmx4k1dNI5Cbz7AEL93eBfKwpTmWbE988EQkMYX8c15HWIdMK
kWNZjft3nDVtauY+Rsvd60Up3Kf6Z/Gh5M0T5FhlJthhdlqYlzpPXCidQ3PLM6aOLTyQXpclotlb
e5cB5nZriRZ5upz/kTF+p7+alVAvuhgmzHHUYlkv3QwusHYDHDcfMUf+2BlPd6gEnb3Enw3h4Pkn
D8caWR0saIwYzSIMpO/NLimPxnMWVYJ10YjtMKd6/CJDT+w79iMfHYFP+jj5xoa8nDAwEJCMAyY0
TNF9MOZtlxO9UcbYWUhnBrl8pP/i+iR6GS/+gO3f3EsmNNmwspZQ3MURW3s4TqIAtsupl0SiNcOh
zu4LQQKNr0Te4O7QX9Mz8doK/GccE3nM2SrqZP5NgCHvoct8T69xccoWI6U4CgzTvel9+c4zQjE3
+oeM0jGys8F5DBy4Za1Km0Zx5NukuCXTi/T/M8I1xSixTHM+0U6Bgpe3J6Mhkk8rCu9T7T7buWqi
YFvrmtaC3zeA8rHA5358nzCe6LTIVTFN8da9AhcVWitl9dc47zPjHWVIVS6M4t6F73SjTMvWdQAY
dcDkLoE+0iSwqkXt9THP4LofguLZ0YIZVGPQuNULNWERtTUNInruqmpLnIaCfrHV8ZM5bue3na3F
aJCBwKjSQgHiSG5Xwm1qpY88+elrwPbXJxidW8+nJrzkATTH63UhZwqT9wTVbg69DDZHePzLUEr+
K17Gy6rnh0RAtNDBEaNbaQbtlLSagwsKgdIntOtM028AeyNGtyJGBQr8Ns6xrqu+e+Sm6ibGJm/e
LUTi8Tl3Gydy9av97neo5WjGXsyQvQJEzOgyE9R2+bYPR+cogLWi4bYKhCeGsaa/h6Jx9btEomEl
WP6j0asAYyvNQjk23y1NLLlTg+PSmystp2cWc7vOgk4v/rqtV0OfNKc/Bqk9jlLPBHJ/80OXPau6
uxx860juf0mJo2TPPkTeOmzzNWjlMCLBR6GmIfsP0mGXbntxlIVp1qNju6bXKHl0mPDHjgKrGwY+
gpCUmDgeCvd4MNtzHg9VyXlRSAUPpzmAoE2AOdtiwnCZHxoUXmbd7KpREb759wvvugq8hYz52i6W
EynF22/Jtv66i7pxkH86SQjYcI/wpfw0ziv9JOadSXzovEhyUtNqeepHJwJ8PtzJXJnFMKMcU9oL
1JLlnjSKWUM3K258Q85LU/BjhGLteOva1bAAK9N7pmX9tmTFwCmQQxyEKZhqhZY3lh4l48nOexzp
GMT5MTlWAeehzp4rxhusEB/B+PvPfAsuRGpZtXlZaAYnn1VGam+XrpF/CQJGVCrGIfzyVqXBC8Y6
n8lpgo3Uci3RUoHJ6/NtoMmpS8oFWS1vwBWyqR67YqqbD4hatl4LY8tNhz9TQ7B8LvXgZXKk5rZZ
brP5v5VncNcbkpfWPtbEpFjh+2bf2Nfm8M9Uqpyti4pEYVFx4SBZSyoaKlZI0tLbZfgQzokqzb3B
4paj21oqY2H5ujOQPqpJqUJPfOD6Y0s/o71gX5uDIvwoOq+xnU6pAL+v4IK6nsIYzJt6LJieERlD
X7BhD7sGhKhz2FOskJ/PJowpiedBkPJFYVJ3KwKupa7XPkVmAByIhm969rMcUW35UPR+9zF9f/v/
xUjbYo4NdvipeM3Z+TRWqhma3SmrB4MZ09pIsTnbw9cThw305BkJztiuCSSnheJ8YfM+EkZO8sNy
G5OIW4MUC4KPp9mQKL2wQ62kUh2NOFtCIyC1DwvbOpGMJqOfwJ8YYXAgCpus07sMXxoIM8bHIusQ
8vjPlN2mDiOWqBeV0bOZnpbjtyv2d06yN9/6Nv8jPfTD59WXdW3HvpHvpjTA5sL/q4HmJvt9jTWV
kUPevlyKOeDqGa+o6gVxpKWG2BnqP1mA4icxg8HGPqhU4RRX4yEbn003pP0qBi/BH51Er32jku4N
wjbqMn4q1nE8vL4iD941pkcDGIqKWRd3d7PqVbrhh82dbptH5IJfpLvL5e3YUecdd8GrIMNAjPPy
U8V1umx7daS/NxePWXd6WTcN9os76ItYuwSUeznCFxbJTJ6x9ZX41zY2oOLijzZMvWBmGB5A2ccx
rwHRWj/FN5cAMApD3Ns56gdHPyZnIxV84HxzUr8EnXxwkIsNCRsdjtyYv5NjL4b83vmmDEF6YkI1
skrJm8BPDmwiVokAMkbpYlnTgxcdVVwYEcN6u2n3P6A/uPehraOalikxvSuSUSij/d7TRAvsKemv
tQZa1O369w4O9ztlqrkRSffXm7tZV6N2ShZRWaLZ4uSE5Uydl2pxLbA0c3v2Q6o9wyTqotXI9kXW
XvxOE72ek/LsyrTYvPuRluNGoUw6GiLjmy4d4UK5f6ydQ1DcxvY5BF8YKZkVVQxg+NRvpuAov+wE
V4nFyhENgg7G1Z0YifsFpzvyjEcsuzZxf/9twwix7j2omuFC65qeRiD4/u7cY7h+eikFEWoc9yPx
lAaxH9uNlYjB1noAj7S3qFy0qOk40usqvom+/xSj9SxBhBwEW/pzaEj/yYQUGMVUElJ+sTXFop9e
xL/bcXLgIbbyyAAjQHRVmgOGz030SBhK98gdIjlMwnXArUkyPdDNUYQFYaG3xGGh5jmXNVZCVZbu
Pfs+k5nIbf2ER67Hv2PF7aRzcnZsL4j6R6tGxybNaRzXEjeBTqJg83uCuFD6sCsfjW1G3z+UIbmH
P0ApJ/T7PjWWsg4urjhxChW9iQh/6QlOYQ+m56UPF/V5KaS0RqmMrgUZwdTe0/rEHoDogFvO9eoi
gCCa/tCF+TRWbH1TCsJusafQFr6PAXDkQT+NtzsHVWj/W7wiNFXbTH+Hu7qmxxDB7ewjjSZ/52+q
Ok5IJvqYZJpwtRDXCNdAGBW9oVBJZAdpkyt9CIAcp8Q+X1Ihm3t3HbdMJ+YESmH5CutjhSflNR4z
Fz4gAeKCLox+mAgjd2PGLC6rAIzx3GD/FHYfjQDTijo0/grUogUB2I3/D2UYBsDItdKHghiHarrd
5/L78HtWq+VaVfMaIj9WGLt7ZAxi22dbSAQqzSkPPeOhAEadjh6DorT+9DKqdXrWhAt1XgCzedry
X5FqUTCWPv6ecMKQ0pl2tbZLRqx5n/9YcTROi52tjkYoIJvj4x21z2TWCmuSd+24GXRhPB9JgFry
1Jd5WhbOdj9TfZTAzzHB0Jc38vh8rPjND8aZ2PqFBuDZUKOXFglcmjawN06xrhY9F3mO7YjiKh5e
eulQWo5rJM5mUobxy+hCMqjRzhCpBAJx9+hguZEsXMGH2iNflAhbpQQE/H8IRTCwF7WeyjmHlifm
Ivm8jcgW1B/pQxEtz5Y9aRqRtPx+fbIGGpcDKnpo7aJm1tYCO0pyshs6lkob/9x0JoJux74V4Kay
C2r/vgiJIvvqn0Ik20UiWvSgXMaSkC4B42PR93og82Dt9JWMr71ErspabVzGlKcYWYJwtl+zIUDp
FDenjI3OPR1CJffXPBT+t2B32rypVb5OhOpRDztNSKtX/BGxPXwXn9vnXvXvfLIJYKMqz3suNoVZ
CBWm7SA9GSMOuRH7O5GxHIPV+/BJFMkDmvTL4nRq8PquKqSRVJpoNRbiK9WyMNB5JLuBkdh1QIkz
/NFxgws2Wk5s/6IXUo1jonR0CGBiZy05pKAU1uoWcjEPQcWBcP9DfC/mG/PYZPmUL4rXefVuPfpB
nBEh9Y23rylZkyOieu5rSvrrgycmnD2t81dSeSbPewD0BJl0EUkGwwKcE2+PhTQlpKwU6eqaSUxa
wWVrUuAey9MfmOvJz9kxoTbtr7v3wA4PCQFLxDYwQsckqF3NuGc9ox42hSCOxlI742NnKzApEyr/
7WAv0aKyOnO0boGDoUzYdk3dzFhKX2P8tFkYfVH/TpMmj4wNUTqQvA+C6QzTVV5sBsquJf0FqBA/
rFCQvBTa1iAdFPwYtqKCe3PvK/3yRbjoIldD4BzhrHoucfkUsWPbKxbxN0zktjk1Iw84vOpiCjcl
OvQZgpbJEGKknezW2+wrgTW5Ily99RHsvH+Fp2oAa8A4mf6u75Z0aVTlROK0dP1GUQrKXXyU2l5z
TisKt1b6ZRBAo9sapHsZmfIiFW1o16mPik27+ITsMpbZOT4w7c/zonDVgWofVyGlMkViWNKj4x8t
Q9JoT86MWAQpNWVg+mS1kSDIuHW7/vYL1e1PRuqnQAPqaTsnnfKY4QNaHgPCSH+k9KS8C/LSRHtH
FMyRivhTwKk6qiMyU35K4n+WkmTsjazvs/Vywk02tgHSCF/v0wYdJVti8lBZ3VMA1sSDrljbZg94
0E70GFQZoqrf27TUyv1jHE+pCAvXWla+Jh5RX1mxO1lWSgtQoqAfTbUbYTLpdy8qjLa5mrM9GYcV
PRTOX2eFjVLHJ3rAsSVFjH6AcfjoqoVgAnUGwRCycuMinXCOUqSIll2xM/l5UBQX0WVLCWHddXut
grUbyEAzShyPndzA/tAXyNBOzKa+ypZGJAXeWInX7xXsZ5DfXGtxtgcYzRTNnh4y/iNF3toUDB9l
jDD6L/DqobTfxxUKNuDzxaJTAwSOY7GG6v5MojLMTQ+d99pzl4qjLQSm6gn+yJ9fd/zqwaM2uLUb
rhfDlnStr2+rx9X0O44EdbWJ9vxBsG2zVtvDtJDW/UDtpqj7Cj2nxqa2YdDVDRI1jdig0a2BStm8
hWDZe2xr+SkTDqbsAfSRCl7a4KDfSSbvgzBWSnc2Xr5GJxkPrWnh2T/S06K9JsjaLhhUqVSWxBoq
l0vZUqNpUIfcaVIlGOuxNBiuM4zZJdVxstXwF8+jwKLCYZehthl7K08udSJhD6+3Ij2lj2eDBr9E
fKzuynl0Yk7hh/5xJRoDyW90GJGPCbR4z7Gi28KlyxEUDljNhM5HNPsAx9d+bssgRBfPJeQP5YSz
p9rFXoR4a4upKecG7soAzZchb1xoyRpDwUgW0RfLXiruubDycOGcED85aAgtdZLc4wqlDGM9qZK0
0+bu59tmxHdnu13T64S3+7CJsE2t+L6ffRINeuudngNbtCX2Fcwo/ffc7Ozqbk0wIcEeli0Iaza+
2V/kaU8FLVwUEje2szXaiiLDFNamyfqIROurNeZCO59pWB/NQF+FXSisTQV1Nx5UsJUeSHxg+GOS
ONWInK5oL2VtWwQcnLKjcdOvYCskyy63VPUfmszIafBMmRkKTDnUr354WFfyRpGpiyuu0Eg9aP1S
a93vnrQMM22ZG0c+MdiWiPpLnoy1m4VYXBDmGdwGYxfodtGcTCPaHSgQlkWCVn8Bxis8LJd/W6et
JXQFow8dvK1zBqsu/v7kp77cMji7jrX2Nziw6QEsEquUdde6z/hol5tLqHpl1jDIikCwkJJ/fAs/
wM9jsYojXX+yh8G+bCcwaOkf24QqckUzU8R5q4EGyYhC2qL016d++H1PZQo5TrMa5sHjC1q3KZ1x
Xw8IsUw5WQ69Yb603tf1qb2YgG03nP/WtekrINrGjvkL5SswthhEYuhIUrXzM+cnBqXsoGh04Mwa
MVmhnGQXON3Q7tlIhvraw1SSg5Rj+isYUt1pxnJjDivXmPeJIKvPmbNvI7dSve4vyzc2dstHQMFG
KiJwzf/0wWSbZJs5/jRav9xifK5PpnSia1uc49gXW7gjSOAAEuUOjrhD19R8yaL0oJj+dtN3tE5H
kByCtXFn9iJm/7ZrU449xt1jyc9rtGM/f4oPkcpZM76wlATaYj2bjJkg9+2+oL8cHPLlmyPMetuP
idtnrBZPTVMIWhU+dhka7a8iMqqBd2x4pK2acIQBWHuH5jmGmVyed1uGFCVCIwCgGJEPa1pVHThh
pgkPEfDzJpWmdBjq0fGQuHskyVyhhahtOKmXnER91vZv76y8cTTVEMRyLZlWMdMHbmPIv9v/nqC/
0NzmQpWF//6cdVovTYNOjkzBKrvvoYYjpMx1TKIDz6B9HoSVPC2V2+nNAJjprkiagGy+GIa7sgur
qSbxc/cjUIlN8E6SN89A8h5L5lFyVKtHvf9lyG0zngoezACxou8pzHqDe191/UadVfoSTn5KMNDd
bU55PBlO2pOME/YbVCA0DgzT8nWXh8qXhk0jH9GIpCXQFp7QCKP4hKWl00Q9NWo940s8bcgQh0Sg
fP1o37QF/a94WNki8dE5Ic1mWwcHe+C09+iLA0dIIfyHwn/v/jFIAYMYI3BnGmkQUA3K4YcijaB9
7mE7SmyEKQAHKqx9qsmtFN4O+4/dKXXEoVw8eim3kD05kqwO2NVirirvTkTF9gRMCzhn5L0w/Nmm
wkk/d5rJNTEy2QxgHSikgqoIhGlRMKfXzAZ34pm87Fr7Nu8x3fhAp9aUSl9PDmWVqfHDWo1Eh+Fi
iIzo2BNKoM4nhoDsbS5PSjFL7MkgFBEUSVDpPmhZ4Vdzx6PlHV9zcQ8aO27TulK+H46hXEM32IbP
f+dEfokcFOn5c4ZfNW7lBtKh0CMubAOFiQUOysgDhcyOUP618tf6GVSQA75VDDelBJkgCptDu89P
7rxpcCQpm3bMvyxi7CNX61ykU27MeY3CWZNHpTfEp/+NBdsi3aUAve1dt/LN3Scy+vPg3AmKOU3O
Fz9s5nhsKfIC8Sx1whc+8ziKlIhok9frbYd3MXLIwCNxFFWLy9Ca7rgMvR2OVxuqI7hsWRxZDtBp
OkhljzpxvwfQWZ3vkxrKm6DShxZqFF0vPiGx8bcNqHRSh40BrKJ9KAU+UXvSzo9WVwH/T+x8Mc5Q
yyOIn0o0ZyhRCal1DiCQSFDGb38hwBxK4NXdCe+cKFZpn/YlZfPnl5Rh8V/a5AZqLbLpnB18ptJS
d67CAhp5cjKYHjbgGYM02IsPA2JQck0B0PpqwgP0MWUGXijwvTjzRj2SerO+n+e25zIDesSNeNJl
acDtizEM7ZUAOCRJNROUOXXby2Tqm5bDd8bu2AkKmHeQK3derttozQ6dJJaFPguLDwFd/X49Nbmo
aX7XEIGYtl+Wuo65Y6bDDSYKo5uDQfYClJLSgJocYPQgk45ufXxbR3EyEVxqO/4EfSLYjGhLxU0m
9JzENNKwcFa3sgyiezf1nw+f0YKA0sCBlAQ+HqZlixFaYRBw8M4GWLe2cKjF1RXUAnPq83qxI7P2
X51Do18S54IfkZI3CQ0+dJQfr77pvQOt8TNErHOCric2kOfwEnSrrRUg7EdZJt3VSp530TSqLXZ0
coZWCi1hMqRkzAGIUCHV0aw7aPXQ4rXaOoBRNeKMJKpMQzlMXmNxbRrOIpGQgJoR8z3YnW42Dli1
5LsnOIuOCJMQO1GmnwwgFRg8zJUyizsFVsjvyJ65+G9HaZuvDbvPm89B7KjWXrstHNsz+v9K1nMO
II+7nCazflGD5o16mtle1wRJDbYM82w1pp34TqqKby0MTYGuNswhc94Jg1x29cUxh9if5n7/bv91
yAznUe4Q/TIYzqAVB7hADlI1uHII3rzRmFr0J74IxPmS4tAl6+vdSDtbCOU9U5Lvb0znq1x1dPdo
9XU1PVZDN8gga8bHDa1tD5sstaGyvwhVtrS9hcZT+IHKqLSsbldPmRaFGkc8nlkNgNZHvvZ0nJAN
MU4olHyQSK7LY9jYy7WQ8aH+aD43UOA7Btiobp2nuFq+pZu2uc2NRt65BYk2VaXyBK7Zb7s8Cx3g
ejuBKhoolzRd1PRU7D4tp1kCxFl4jM+dBUPZv3O9fa1ZaTKjhVbrqzTl5Q9WoZzKwti/0liE74nv
4753VXgTe/TfWBfYhrRZcllPHwuS8AHAL1f6iXOqSEhKAUqlBHCynHpxaGJzJL+HJvmfD6Wk1Bqp
1tqBaAzRBqP/TsYffwlBLfqlkZOM2LqT8inLBtKBtRJldumGSBAc312Vypl2xR3b4zlg0DygjOBr
Te9G9vDQOM0k8DVcYuuhmbs0ldwAljelqph9nt2MCdhb0cCZ3WLY947Mwvgi/yaxDhuS2A8nW6Me
EHQpidkNTN7K87LCZPiTjRDiSlsdIRAvqwWOmrd9vHBMAD63vKWkyh7hiZLXH4skRIaQMTBq267L
mYgQD1SWWQMQh6dLpVTQzqspt2g4XVzk/fTYtV5Uwvf5oHAamxq1TjOwLUFCjFZ3IouoTniNHM5k
1uUOvr7TpHaHXpszi5TkCu7GJlOMpQg0Pf6k4p3dcbZhpbEHKRrRkSG/rpsMKS4P/5UQJGiQAHfF
5SlxPWQSbwxmX2ouSHzRMODv2+0/YFdecLSCt6hjOJSFIchJHZziwhHeBi4ckgB9IxD9L8nVILQg
/YQx3jNWiupPKQCDvrcGQaRs9eOa+amSFH4StQPHoS5pQpMVZa7h0UnmOQ1ca4fwnoTBDAX5VrTQ
sxb5xjacb80XQbtKx3FbmC9ox6EpK4AJLzRJcHEO/o2SAFyUiv9PEI1yrzCInzJPrTetFnwyG9dN
ruB/PjFXPqtlTyC6pIJf0kFRiQ12WN7YaX+WgWHhQzx5quUnRb50WAupu4YPCV5IYpf4B9byxR8x
vDzZAKIkeczFwWHi9VMs+TFNgqWYZg2jiTNglrF2XieIHFnmPdwhlWW0bj1wy/JV0dD4M7tGLT2c
6dk2ekUPMKpO2PjOLrhraLf5rQu9V3mIj5byjALSZcqtseH4hNmuvb6bRB+CPvCdiSWIKZaCkld6
u99+Sopvse7ZNGdQBq07iHCPOjc9nG7Lv2E4DS+vyPJrtDjpgnr6jkYQkkTfD1TsrQtKoYHMpQyP
YciZpyWuP3GdWP0xLxjIqKG6Dk20HAkyOX25Z/r6BTWB0/r27f4yyO02dn92aMhlPDJ6+UiUPPLG
QhQEinBi4GyZ4fDjT9Q62QhODAHGl31suiFujEp7r54UtBkDkWIQmE+Pel/R3SnLeEhA8PByi43p
vdVAHMoXnkWdEZiroTWjE62wYzERE7SfaLeSyK+1s82/Rg4scOaGI2QTTHjK2z77FDiiWcuB7rqR
XIvQaA0grUdosmiNxC4u6UXdvTgSTEtEf9A7r91/csXIlEa+Z/DMWOjyIjosgc5px8/yinWay437
AagvIYBI7Iz31LSy4kZ51NiTV61hJOPupGe4mXzVm9xwNtDDYbiiH/7h25TJGZbmbM8i2f3Gx+fi
MvUStrSdCZ/jqghwR9286NNzAc4+vKR4MBbiu9KX4JeEp3tZB93/BohKlq2A/ZnSa4Rb3UMdqQFQ
khkytkzPxCRTHbJLlGbRpBFFLCgRvXobYVngOidyj/Pp8Tj3/NiEPopibHEcm3YTv+01BMxM6TTh
xRwrYk4RfBdpEcaHQ+lkIH2ycEJ/lhOgI2W3flGkauiP6xRH+md/WhXp9VttWviCIOoJUS+D+6i8
1ZN0uqONzQdyt4j4mLUlW8WYq6kK8PZiYK5MQNRtq0vuvSLpdozvHz5QBr/W9/Lb8n7PYqAZ6GYG
P4AnAXfcw81GqwEU9XPLzJW2Ab8U3gFuIfpfwqGqONQ2b2nJAAbzKEZvvV/3lzR5UTJakRDkZ3L8
WpucXq4Y5EF7ZdEZvVfzic7LlLyJY1571CvmPfL57cdPz/eaVYQ5uPfs2FRjc2mvh8hF/eVbXPUZ
0R/4vr/zhRqvzmzhIz6iJzjLn7EHgZrBp8ru+9wnCRX+AhnhVeyU+aNVXIZFQIgJfUqH7NZn5tlu
efxxZ5BTsbY4X4XyFPOhrIsB/o+uMbuIwK1iCOkuUpg6KeHu7Idf5vc60oKgQ09ia0474fZHci1E
P8i/oc3CJ/K8m1e7fxu+ho+YMRN+L9f9Hu3Z/HN72FBGsXC85bTridB4owQOF0KqNVyWaXSgB+VN
tF/4YcsqJINXjVSyCfteMCCopB+3JMJi5SIZhsoO0KH2vPZvvGRUT7Y4VoF8GWOMKC5tUlRO4+xo
9Nu3hf3ZCJZsiakwtbMygcW+DKXgU6REYl+VgFkpyFrXvJBypL1WALeZkTmGlmlvC0buRkIqUb5a
9T0PL0em+T14539ZBac34+MOHUCJXUOTglRVl41FTaIZnCsF3hsClJgw18cCvEMqsHLt7OnRxNGI
B5IorMT3TT0PwK7Lp6MGe9PbanZuphr2iJNMyYiD4dFLSrba/XQ6isakuHb3+KAUqEyVFG7F9MNx
9WOx+84Eigpm9zj3DxTlkbMqxRKeJHqf+YuCLT/IEgPyvC7bc8gQkcDF/dFUIN3NnmJe5F8liIGV
hmx3X8XuaBIWz5hnIGE94R6+pI+thljEvx59xaKxiztEJPxWsLUFge/8XZNS/AOJYzdIm1CB/BnP
0lGNf/dsoqZk2S6SexB+vNyvUqzcRW1yV+5ESmI20aDWS3AaG9g29AoD0sU05Uk/gjc+v6T1wJIl
sUogcEzTHJS+llbDizNdSWbFrwxiOfinpk++fxJWEiTcqBlepUQhvEoXFq0yMISsxXF7ZWH2dm1w
2GCtxNK2Zx8IZEMHJ9eL/KQo1pTvOPL/Dq4aLQDC818PRHmNW16AiKrd3EJkQ2nzx2qDOsUYH6w6
Wphyqlf9qcGi66Ow5R5OiNSgrf+T2EFJSKGfpKsvt3W61Lc6TzQIq71d31NWhUvvlOYo7daflaQk
BAM7hKBLALdieS5eN6BF7rtBb6Bblej7lFYV2Jm4SIATGVfmVyfynjw8UPzmNSskIDj3LES7TmH1
ITbXODkbzbDcjGgHrDlmH8uJDPQo4U2Knn4/oaqprCHMvx18W8hTF1HUUSrfRtGrc3wuINqGoREj
7NKl8Om80MsqzzxcFTxPcYEyqI/iF64ohjle5A/HWigPuH9Qk/Kk2Skxr7b2S5qkDhnSX2XKH1Iz
cBR1lsiHYF2O8rwLWTmfuIHrWNsMGJAF7lA2GKBPaYVlI/T/dwkKNX55BjqqHlTPcMHxbOnL4NjR
hGnagtKsSfcsYkJiiUiXBLQ/O9qf+r2V6jLBPSC8lkzANprLvM7zemdohvi47f0txfydd7UysNaR
miMVZ1Hdu9Y6xEjoPhGaAr3W/1XsG6pKODE2k2PmvVpEqewzrCqPeu3cn7gikyEuQv0JscIBa5AM
RxpYj817Q2YPkuZK5o2nubnjH78ixjqKJwEFRjJViU5x3aaQB3qqQrETZlaNYXBOoCR7/RWZbLtm
xT0vMNCV5DVTVXye+xUzMgiYrVL1Fm5Yiw9WuvgLF1amIvscCasIz3qMPjAE9+WVFs0GmOrrDnoz
9d4YECcWtvlPKrqeN0Z97m7eXDZBKlVvZdIZlaBXQaGpOfPBm7VLoGLoZnjMXFS0SeLIvNaVc10F
p7N94WyIAEseFTERKoivKgdIxePEwNU9PbUbscNf/9pmpV7Mkv74rL8GlnbwKkNu7+YGo5njfAib
paO8F4UT9BcU4D0FGXyMi8PBxwoXelCR22yeC7YTqJ9xbvMQs1XRVpe0GhNXOk3f7YWq8xiHeF9y
5XBdyO99vbkG3EF0VhJO4PtMHFK0cm4L3IVyhbnr6b8VHXbvFBOPIlKHoDV8qVMWdRdrcmkNhbcX
T8ZbtsAJOcSE3tStZePCp8+mkcxy4stTW7K7QhNzoO6XFuB8DopGc2i0ymaBI4syqGhYlWcVYOn6
fYopTo/fG2ewpV0eSKQoQOVGpTkhVK+8g3Ethu1VPVl9PDYMryebQR5w7ihKEUlrOM/wVZ3GgK4/
68Gssf3h8p33ZcI5+lSD/GnuLXLTM/oI4lF579djTVQCt5lb2cC5cyaGI/aC6iKhj4yNpM8w+WB6
GheBemqtax6BP3w901CcZu0IIS/PstLDMoG8NRtS36ApTWfGluC5MW61e1v4gqaGcCHNlm492lXv
vahfR7FylmSSt5suAZNCRsf+U6s/TIYSjFJ5KCsnoJn9vMCL1Ko0pbdyUlQUpd6u9BtoCwCytqQc
h3dtUVLeXwBwk7nnz0XEiVwrPqiX/tttNYjwEZL/Vp9vq9tybOXrbeyE9zADeqjYYPZsz37kJAYt
ad1tUve9+XJsoIibvIJIdhQAFpgQkX3u8vIG09bxjtH0lvpjLy2UZkgf6qPq/YIimnXpynQ52JyG
OdW5Q6ninrg87F9TNVDcQW17UoFYEl/pnF7n8OtewGDBEgskTC5Wm+ZSvjALGFx9L8kbGWpmZ7s9
PK1qxa9+LCN8m3no/egsWNtILaoDyB9ihuAzeS695MX3xLUdWsMGyC2uQgzOtMXDXz113sbN3EpL
+Ypth5WZQLTj+xubs3B05AoN4S9i1w+RRWwtbIGYKi6K5zPa6IGVhZvnoxcdrISrTK5q1ZGUJnVr
PFcBExABkcRMNvU0M8adfHQx7zpK+LX1PYxxo4iHZL26Rbk7fx+Rygi5LqQbzUF0vxXZu2yW2RXC
wXi+AA2dB9CSAmjveR+lRGZ2E9z+vmk9pCFygxYQB+AiiO4TQgM4V9YFqksoLwL9w10UM7GU5Nzw
6aSOv5gfCKC/HO4myn3jFFcohEGoFX3qL8AHcFvvzhgFCJuw2t7K4atcPlb3y7e2ZgFJauqUhLan
YioyM8f2Ro40bPokEBpmgHv7uiOZjkCXAD05IuWW+kx8v/Y8A1JdbxGdZ+UXIDoQnUX/knjfmr8g
zzbhTN3wHlU8ZmmWfQ3Q6icbimanx4WVL6dXAMrJdEF/Fq8+0OY6dzu+Y55HkU8pnTREU2zw/B7F
tcGIzDdYsp7GdBHpZncljraS0Y0UB9euH4HShqsYThXH8BE2IRPf7TcrvITz7NXJxrdiJCORWvzL
7l69eRZMQmtWAlGGE8EvVBHLe226vlUtALWow8VJaNraskPbRjvY87H6+ezowFQ6PM4kQWMR4u1i
9tLlBJGd8St5F+6Bk9/9ax5STPFe/KGq30OYNU2fXn4rTGpXzB6M3szf+PSniFSAudYM9UYzS6/N
92CsSNvGQYTFXAqlHwK+w+QiEaKFgm3HAkaTpMG3MZpP/bTP7D/TUqkWSjo3pUKijcQ/RoCOK2qN
nt23mVlo5Y5zi5vfhJylzMG0EuhBBvxyJDQITAU0y6SsXPNL8Wj/I6lqLb8Ymm6WJF73tDQDkHif
INjJhR8uxhWb1yYDk+W9y9VglPzUKVtl3QQk8kr8IpbS6soZZ5MEs/uPqflz5dfVceWB5RLm0q5e
5m2BbOx84DcDKDrB9mSKD+IhRdtOBC6VkwtEji7XJjse1KWbcyLsH2shdCL4klnMAqaeEvTaQwv1
yCzIT665kMYqekpc3ImnOug2t5Avg6aM3ZFasZg1NfXbrqVlnSHPTA0woxofcSYPKue5kpife5P3
L+qYZ/ZdpWhA9ssV6tg1kRa1U56ZmsZXkDEcaXP27WimQVPpo9N1zSFtF2OMJsR6KP/OGhHG53se
SopPCG1Uas10X8ptq87RNGcVI4vbvxlPbxiXYj1Qj2jMtLkHO+iszuDA7XRn0ocklk81Y4jdYcLM
TXESqcfQLC4Lu7NPvQKeOMaBvYtIeDuEXw2NRWHU56em1MtimUX5fB6qE+r+EODsjBUxEEo1LDV9
puTzDIlG6R0dHtfV5uw8mLoj3Wbko1DhY8w/0eT/Z4FyJ+tEPufWsZw/ul/0ZT1rysuP21p3V+8J
pZV+73oCwCz25AhWaVY8JxMWq+dQXlx0rNYDqjDMX0nrlrSxSqeTJhyYB9UJt+qqjZ4ExXzQ2nBo
HvSPUxw8K6Evc8bc0GSaYEUApUj6Hoe/H2DxZ38Nf4hhnB8lqOn3LCt55kyFDK3AnuirzMB6qHbx
IwmYcTVOi3GfTIf/zHFjAkAk4xfC7OmJpUy4R1Pchm59rjA1BDhl84wo6eKXGJKLTmYlHFGaz6UJ
V/Ff4Uo39q41jhmz96Tlm5RnMpDB1BkLYK4VP3MGG48DdoO28GYcNuX0k0WypB24THxTzwu2cGxD
wCyIKzLv3JtxceDr+MhaDZ74Pr1M/xUtOc3qmvC4X2df1wvJ91YUP2QRsrxqtWDuSTrZxe5A736G
OINLF0drS4hGNludLawmZuf14Mf6EnepY3C7RbdtWHEzrA03UexIxTH64sseoM7WV7wMJA6dhkV2
wbnE4lwmMnJMxBg/y9pJtfxM1xPzdwPlqUOSbRnN3TQYvuHzkVpPCmiNLcNVWGQY4DpppH7eKP1F
+VKItlzLwAtWkWx8osebsPvfDrXeG8uyq1AU54K0ISPAteGWUBnzQPl8YroQPHizjQpksAWgPvm7
t3ERAyqPZLHieLQbRU0vq/q5r6hP7m+OC0uAoLz3lbURcscPSsnHrwtLpyts9Eg/4Zf7msSyDxUU
nDd2ng6CBWJQV04rDOiwRJHcgJ3wJOGegBYWF+LYBTjFpabqGedP+vPFlCZl3bwUesT7/c1zCEz+
9NLlKL69p6DrAjo/rR5BDn2MzY40v65grJ8clAS3CUheBGTbyFA0Xqd0yr3tVo+jPCIykJ2s3Qzb
jdXR5p1MXy0BSOiUmCCtyh49ABszMi7Lnx9N4p17jwacI6CF6JTVRH/mXWaUFpRiJV4FBiTOrCLR
/e7mgB2LcgDmJxu9d+QrSqqQPXF38ZI4ZULJSd9JxfVphffRXhnGsw/cSgJ5DDluz5SGQ01/irQi
ZbQsiRAZ3LQ5F80ioc3qZIWZWuEJ2kgbqB+6BRFH6ioPGAnbQf6FyBzhRtN8qjW7+SN02nGuHxPa
HikFf5CpB8wbYfQ/08l6VrFIj5lateow+ofxmBHUJTYSiKEUAnzRncjFdsmqnLk6Ml7LHcIU37Ff
VyTYxLKbwmKnVvcWcT2eu8oHnT8q3sCnA5KUPB5U9fmu9+v2eMkSJ1I44pbWxbJgP22HtlICFa6i
xjznhq9HHaO5WVZ/OaUSO9jYSZN+fbyd6f74+5x6w0kkDFO/l1vvW8KpWdaVToj7pK2j7vUqkMwL
WinTVfQwgM2JTehPMuVAb2YK66eWApb9qYTOsHcSySto6q3YcBXDpiO2M4hu8rw1G1CJbFHOoWOz
EEI8Atq4sbE5tEjhri0vTT4JixaZQiFI7+uGAadHWnNgdEPBxXjIhBwkpQCILf4Owcuetf/UiCMg
W/tvbJoHncf+XKtaWSBlHZtOqM56rbbV+uZTQYA0owRk4f4paLWcG3q/659oMy+vBVIIrE3IEfKq
9XN2wlteJ0M5tDYcCSvWJF2siwC4TpLdd0gph/E8syp8UAvFqxkwWP+6p5AtyWRAcdgwiXrrKTvY
14rsHByAeO6/bTReB14YmAeqYVZFYXUDVjpmbHpPbct5LPOMJG+LyIJdaU7P78mGsU/W4eU8NVSY
XelPZBlvhISzz7uJIjF5Au5oVjCvRCrHtLNOCExy7zHgu2chx4eYE5sJzDVAW0aeTpFf4eQ8Y+Fa
xz1xZ1pDITVnIrAKiY8Hh7PhVsouiO9YSdXl9u+RxSL6Hd45uBf14tAUOl8U3kyn+WEslbfvPKog
ldUIMmEhBk0/c4DQB+QDFhqDsYveDWcMhawdoerXWMdaQHNJDd6Y91mRLmmNpaobe0uKqxWg3r+G
0lQWxttnQlZ0JrDvdg2W/7Ir4FSY7Gxv/3zOm+MOrwpNGCTf9QHSlih/hjgF/AHe6hzHKdn3klqB
N20WuhrOE1vNLOURlaPO93t82p/UPk2XrVTZx+KxRZTc4ts1uQP38wY5nkPwZXht18vlDImCzcpl
RzJrkZr598FJQayeGFsHrSu4vUdwKnjOY0df36TmMMHP2uW2Ng2SHpFnLO2pJjq6nCNxZS2SXp4K
T4Q2JF67Po4TR9Mt3QqSu7M1f33DM55d4z9cZZQPh7GSHcsPwXudAIdcTK1l7ZGBzlnuXGsBCMEF
FjmlBjkGNE/8M+mOQdWpY4QfrZv0vpbhp34i7/stAWSPNzAtQ4WxIrd1vYUEAd09uPh48Ek+Y+7g
OO4atv5JM+0H9+ScrJisZL3ofmNHjN9jC++ecFPw05/0qmzUlMQLTVrk0NV19/Ihard+eGALHpAA
/bkPGm1T07y1SJ3ZMasp/CpuM3tElk8YagGu1TCfbftE49V/u+d+KcjLhhz5qX0QtdQmVW1UCeHE
ymIxHFaigWZqDixG04IOQZJvUEYMMIvU8PC2d2BwwTbiOTYlkWf75sk3M/X59UzYzHkodgfvUI++
TRhB0zZ1pOy1x5rljZObZ6h/PUAt9Ipzohqd3OtdL16di2IPSIfnlYigTy0XY0FP/QQKWWDkhDvq
ktEFBDfwkI2FgxcbeIu5EObbOz6ODmHQguBkxd47ucNe0UVm9lGgwD/mw5psF9VE9hF0WSrZP3TM
BcmfbxNy/pUHRZ1N6wlUaqbDyhv4721I8IuZ0BUwHFmHwyKohzK8WlFxBcA1apEulnj3WMxG7Epy
D3IuBGxaSpd7kOJCPCS19rQLStkC6b5n353zB4E2idOdRDZnC2IqS8H5RfiAgAMKQXdnb8HCe6ZJ
z5fOKweqLsUDC0OYbxr4LCO9tFPAgg8Aw/jLSVsK8DW1uOOgI4RG9tr+5VXsp/hLiEZsg29OyByH
pnREWfGMzMmiogEP5QygbV8I65186S81Lh9tVd9QhQnvnTjhDsHxLekTdnetwtrKl6brM38bsvKZ
h5g9k1VbVTyomgmVDP5xLis6xMKYNIh1ICTf2qvit+VJXxliZkZRDn2bZ4vigYUVhvxw2nFVuwJ5
WaDftws4UhGSQWuL55g3vzcrLaAk0IiFJJJDWp9B+EZVVb1J3hBOnDQvRDt0MJFLTh6xGLt0sqnn
5lBDzdoPeFuv8ODgb8cVMzU8wfA/Ccmwxs0vShMsNWrHnNzgaJs1meamFn58XFktVdKE74MUtb+p
VxU0fP8iu03umcdz+dpnHTdwNVPkLQokyA/yaCdCZWgD/EUk++OT5JsVDnPGXfJHzXhWnNr72QQM
n7M6zS/hIldBMWXgSfj3JfsdYpSG0xJgQF8S96Rv0AQ39jxqQ1b9t6wJ1Jl58LH2bnQpZAseFSrW
TORUq5c/EVH3X6suQASeo9Z5kQoJ/pJvU1YAVrYNO3hGA3dImWR6CCLptw1b/3u8i15wNCvoO1wi
OgcAFCwmptGz8PgSfml1ellLw6+YiVeFEU2nnxjlHCQDO+8MwvCiZFReEZMn8tXql4kHTeEuZ3Db
fQ2uUSIldtfygIl3zTpFuXYw2OGNG8SsNFQL8iw93MUUdZW2JNTO6jJveLZQdVY0N3gaAI74fKXC
qQgO2zqVl+Uq7ulN29KPlAtmymYBXq+78lgdMX1/pMKQazsc1Os0ACpg925zi8r+ZAkjQiASvUxC
5tlvpKzg57dVdUCaxqle1ckQrQaaez/9YBUsGO8aALzyyRG9otLRY1aAlYEDmFODewkAc29RJH+g
hx+p6E+2IkAL2szLlgF4xJSNyE1Hd/bwaFCrC9ty6ZJ/GsTELy75vB0acnbU7IZuFzaQ9nnYD+eP
ubd88uWJI2UmNdMeP1PVFjmiz8RDjGNDAJBS63A4BWq39Yk1Vtr04J9BT5jPUYEW3c3hWkJCOVP2
kLn+IPuolLB05HwZpkNEzSApJKEZo0KxQTTYe/dB0TJXBLORvwWToBib16QxvtMEziYSUKctDnkJ
ILb7skXKFt0L2suN46s37k13vu7hv1RUbYjYTSu0/flWCFxbQdLm7QHZwIPB4rMvMyTmOcA5yZiw
xhz97LU07VtKSYVqX8uhSzI+GwwsvAw9hE0oxPGxPLOkfIW7q5zwlg/Wcadh9ZA6SuYrsCSO10Wg
6hm83hWoln/mh1vODYKCRcnq9rlgJbEvOQuJX7mvgBl3spgxRiIa9EQ21Ya3BC6zbB3yyC4bf3DS
IzcK1f+VN0q5f7mJx14W8QTMrtH5A+cVVD/bST6zjDgv/CsO3tZLueAr14Nk3HFZbbrTbgqxbBPM
KaNWEDtTFsgY/U7QLr68Q4gok/ZA0uIdoz0hAnq7Xfly1EXRMFZRRaYyUTszWb9w7vvHReBBd9dC
yjjoiAqNszdBMVfGLFUxOZem7IzUrtkksJ8S0LSN6/db2fu+yT6yIQ8V8HqtsXbLMSecEFxlvs95
NPwYtjxHLHqxf4BUaPOezIUALv+PWmljtMvix5s7DJURIENtgALsJjsoEjvI9decbE7S+QgfACNO
1uEDXz0JmMpPI5dWiCvk4sdpfytg2gP/9fhvdawZkMxCxJMYeDlI+fV/63474dvyD5EP28mE1eik
6kF5nwlvaP3d+3OUW7rfTCXHMTs1QDRm98+ANiENYNC2H5C+acoHrmslJgn5vkjCOY7fnufcSe7F
xaTbA/Wq2Wl9DLBUyGAAatPsOGzKANkJ6Bkqlc1Cjhhq+Re9RGI7EekXULy/VE5je2F7zN1J2C85
QOuL2IqWfAJZcRAegiMtaO8Dz/n7hbEQ/TcnOMe0zNgfwrxTN9+h6PlDZugOGuqhE3pR45SD6uE0
PhksIENtHh8UF9Miov9o+azKxZABEtCcK1Rp/yXQ4u8amb6k6N0mbPNKF0c2nNb6Gx1DCB9ZzwTR
0KpwSPA2P9BHy1tkF3ulOVj1zLw5B3SDMPh+YCWQtbNrMFjszZxheHedJ1v2SvzviRuPSM3e1Xoc
vV30yuMcMwxOvb/Vh6dYbGlCKSTgXd7fJo6Ew0zRwd8cwhh7Z/4fypGn2+s862jfbfO5e8ZyWZXV
qUgX0HJ01L7ywi1CpSaQWV5O5P2zCxQkwvLUWYzjWmbmRSg8sArUTFiDP95HGM5FDyLuqUIdc3Gz
mHXZZ/oeGF+QDeP3kiPZtiho3n0jSdQqCZrRez4HlvpdGbY6UNwPSiDMNUqmkra2g/7qyKmHJrKF
C68YPNh0+7900gaIbahrnpi0aQKXSu8VagxLUQ4eN/PDeDuaa+p1VuHnQryIkCvb+B86dbL/UkQT
FKyQg3WkkAO1tt6F5QmRC0DPv5s5iwr7MyOgqDb6JcixOLVP9qW0QEm/3fBgyWEPq/XwlyXhAqlF
2KYr1upxmkKiEAtpUl6omETJvG17ZA1GQVnYcY5onwinFJDqUSy771TD6uLSVL0QBPFO55YtkBJK
QFgX2ODkk3ANCcYv5NrmbHEDbf9PiyELInzMtqNae4z8xNULKh2lcHJcuvwWBUNHot/Ruf/7oDxm
gNoUAX2weedky7GyAOXhwRoHyWjCROnhAS3c3NOS03rO4WYlRU538oAX/3affz1SsqMx0erZ0CD6
FF9GQrkIo1GNggdulQy7IhJMkuQuOcQ8zOAwXP3YXB1FaddkiL6Nvd36pOzJkzDnMH1ik6TRxgmI
1RtLei9laWTcpsE6RrmFS5Maw5jgYo3cRqzsZlSWeQQw3X7ASg/OKYRFebCDPAhZ0D842IKZQcZE
LIi46NgFKhei3e39wPDBfUkpmBKuMYNSr1Sf8nqWpc7tK9pNDG1m/iIZAmKkzi3DR2GL4dWAoy64
kXBYRKPZSQ0tGiqpWxtbNGuyGjxMTSWLKzCfeuGOPbiGHBnk8xNWG9Yxmw5aUbxzSDQd4g5IFXqJ
8rnBJdERgbftvLROufoCVHjVHSSIsgCQHEv8rL89c2d+twzIyHVya9Z+9c0AvL3N6DI4OulfaNNp
o9sWm0Nj34pMM59+MuBElIduc87vVmMjIA3rS5qnyQcXqfVDv/KDrhxnVEplLyI2C5k7aZeMaoUx
5CCouAd4QsdoNTozOy8rMiaclYY/NZJSpWcrBZUyW+sxtBgH8HVlK51IuZeEu/7ZaXLphKgooHrh
LrWsG30wUzYJYhgyTe61MJHquzp41iXS92fEN1JzSNh6zAgdh40HHK4sfxXwU2N7iczAovZQbjKk
39WzLJEWhTpRxgkZY06JFyznx/7pYwgbSOJqMmg78KPkZgpjpsWtZYOa6kAKmgrS68jf7e7NBeAt
oahn29LvhaoULUJiVbBY99EWGZgYVtWSM6BU+Zr7AuC4qr6ZUyTqKuV+BEhJble5I9iDa7oiVSex
hoF4yzDV6cSlV5STwQRmsZ6sOr6aefDXxJvYZhCT/VY8tIUGiZkDQDKylmn6s/5O7WSkPQZwFDbE
1ulaIsTdxH1ss8oRwlvN/WHgA19xUGDyzPu5fQdg5I95bePXbfgQ0M/p+kz/1QA/kXZ2pSDjZR0q
5krKwliXwfNFvt6bCfSrr80n0Oxt7QA48lUJnnf5OuytiUQo8TYHxWPUKR7GU7j+ADW3X113bnFx
B39ELNEkSabB1Sa96UweOM/RQ4Rsh219M4syrWUaeFSMkz/2epJFMgZgTVFiY+BGQc7Ffi8tlj9n
72rzSKLKE/d/4iGan2zQClI9RggyRgdpB5+5ciyM2Ogq9ejO7jne+AOntpgb1EH5pJthuvbQIZm9
Zozjs5eQmvCL9ocZcLNdAxq6EekRHAT9zhyGyphp1xTHvibaQpmcE+Ye8TJrrH3kLSlN1Ktup9xl
5UsoYPoHbw3w7+xIgZTZ2/sG3Ljk8pkmbTg56vsQA6zVdridfJAR4Eq08iOJjDvt0PpAFsO1AyK0
CgIarKh8OIo641tcEYboT9/mGEb791g1YIiEDy0wwIaeXfzThRYBamP2e+bkmW+Cqm393h+VLdyL
PcsnfhAKkzKF1vSUBDtWLYZyPrIkFw3zpOYVFvnMtfc6DUkxLaMTFP6Whabx9bCWy1XOpsHaQ8Fh
PJE4+H7vXnXBaQc7wQDjvBMGYlOvCKMMYz0dTDHewuLuRras07tfa7cLhBwlmDahSx6jBi+/uoEY
FALPZ2Rm2uZQKWqlVihFoktcZtvrNDp1G3o63ruo5WN72rp+7TX4dqpjauu6WqWCsHtW650/I5gv
sU8BBFscaxpsYdwadYx8qE3P+3TSk032OeLm+S2SjWZEmkKAy2k/qPNcDsPu7SriCeksC7Knk095
pzbWrasPT8Ss3Zan2a9cZTnUhPN3MUV6nf8Wh8ybAN7XgTa796n9fEauc9sBrrayyQQtsew6g6+w
erL4/tcCzQfW5Qlm1/KTF7RF+QbO5epixPoHC7eOZZLw+oCov8dQeKoi72jWOmlyc9Ju91VKdQNN
moqB4rNWTItxRCPviqGBoyPlraHgTS3meRjvAl2TGwkUNURJrmvqP6dzwBOSAXd5Wa0C1L3XantK
irVIMoAovC5ODCZ+tU8DjeeQEOKK4th7stgLcB0ARE+gCH5rIbrEDYA1eIVQlUqmHK+GKnPPSF7a
ZLzFb+P+z6swjnyvzCj1SZJ1DrBjkc8BIc1Zm2XRWSrmulZLaaZo2bTHEpo8vGuo5tgLeGmeiHNZ
hMikdI/NEaKu2x/QTfsqbXxeapfn8jI90E2X7OS4FYraHk3YPSZcEjOq9YXbloFi3efuSUTjVkVI
kdXe6ak18toxeQTOUirkPI0KdCjytwzKUtl3lcCPVKtCKwnDArsz95FYTFbyOrKqRsMYjaBbu55g
uP++ilLvsFOP9DtL3lMGEHA7B+BMGr2kHXbqd22I5Pw614iRTpaJHqJJdMKAUOeD27/8E13e+HJr
m3DoF2gHyJ8k25vPIFssksTNIzkqIV7kB8HsoXmpo74I2IFBPff8N8IbRT9YOzdcooDOtcmK9yzD
TfZBjBqRNpM2Aleyuwam9yOKaNT2UPZnxzDh64MF+aMxMXCf3JCke5RcPLfPg+23OcphWJJnc8GO
GqxFslDw8SHK5IrbSIjlWkLDhLa24bEWz9cijc0Sn/U6ck9MJamhtz2T3tAisb/4o8CNvILyxtor
PGjzX/BA+IZ4XPm3laQvh3Uuu+NYlWaz3knLgXpxQid2uHc3w652Bi5qPxZQhVEn2LFVnOihmylF
lan2SU/H14rvtznODH49m+rGZMaA7FxK2vOoBcl+N7vr8Irx58b09OKThIKz2zopIC4LW+9KVAEg
fFfjsY8mdS+BhnCOIQUDgoSoJEl+svD5qSAxhawnsG5/WO6IornFHwqsWnMSFAbg1LAMmkcHqmV7
lkt9H1JJaCstkvwv063t4hVpp7mLmZ7sEHkHGWMdxTH2dfc13VfCGSmLqd58IIx91uZMsWRz9CAO
t8a1i2QWNzM+F0WiszjprzQg/FljraxZ+GotPW1JzYLurF8hdwOR9uShq0OFh57vuRFrau5U3OaA
pMDCA8uQ+Unh6JPQfyxMSpadcGfJeGwfn598p/HQhYo88NJrxTvetZYZ3e1ntpkSJjdC3rFOu+rQ
Rc9/ZmmWhEVO4VFlUf69A/0/Igx0FXrBof/eRNRS74GLqWN3G/zx+LVEdD2zgFFk0Y1XWlB8d0zm
vqQn9myH5Ps0IfcPgFdmF45ekPMHx0Cr3RqYAG9jxBmerChBLw8lwION0yofI4rDDpbsSTfYIkfM
WWgCcP3fdawBmSeZT4xgpwQHaF+kUY+mM9NWqMw0uzFo5LfQidRs7p8Dlyy6jkW4aUQZyX3uTyuO
HgcPIKpb+94gUbMa88WH7rzxkE/cOL54eLjo6H6v0scB34QIbFeygilz9rzt2UI8njmXqxwVHcq3
1+3zbqIANjgvDNFpu6L3zroPXOpt54eWMm5Dyl92CSh4PzIRmduLDxPNN+z1DGzvD//vFmAgIG5R
ubcgI63zXau/smSWkOIEr163fmJmC8bAMN+Iv3PxKRuh2ZWC4tq6q9i3HulJkVcqLp+WNPn8LIsq
4HpTHNtVY3zwIipdWHQLSDye1Wc1d0l4wW81HGt2XhKRg5QcFVv6n3eRJ8ayuaGaFHQvvGRsSK5z
YsAz7oi2eqj0joGSyydve+uux27Qqw0BG/oMk+D6vZUE0KVf5ACRaEA2gcmrCFrKLQ4Uug5IH0Ca
7vvcm+JJqjsQaGs0MXhYHwPBx5P+Ean5q5vmXTmiNJd2kynsq6XKz12W+y5Y+84nj2rq44VDKZIr
u1BiJAw7Iu2aTGOvKmqEq3XG4soNVFudb4RkMbPcFPyelPEIxqsFyAjLa9v7ev2tcnwhjjz5fq6n
gokjPILxaU0HqwAz/5Gcs8B3C0Hme1MexEPHQnEfszKIXNwSNNKgZ2QqAnu5BTRdBpr1ylO7J+b7
q8uXHe+8cp2PhiD8SZd5RIFmDVGyIoq0mhmNzCVp/HOn+/oop8J94+4t6D5udeseIS2UZM5YTupM
RcCAmzrrJv48lwt2r8peAj0KLr3sgurjJJjhjpF5f7gUO4gW6TsOwX2tr7YhXhp1YVhrTtvEn9ZM
SVQVgVQAcEK2Giy7gFGV2ORCf/BKJaUYzJBB2vNViryMguJoTaQ043rRS/boYXSyxrZwPlWkz7DT
uIH/xKata7fAbLlKaIF1ls23Q/AskJyTocg/cASYGsf9c5hoEjQzjkiKnhDwEN7zcy6JXsPkGanQ
LOFELNwiX9JFVTyVJe1S0W9r0CdhOkHlhiVT5477f5AC3QIj62H5fnXMQi/bFBaaU0WbFOB93kGp
vR0qmeXTjcv4SsFjgLximte4EIJGGc9voUWfT5HGM7y1QWkCK41QrFv4ebC16yCTNl0g7rekpVlf
MEi0+bKTYEPuT6X6uhT1yOazqQTw4T1MHDFzFLazDYExrPCQBNeThBlPAZdwxWECIIVaFR5DYyfa
PCrmFydxBmU71IiPFj5CZMakTcgBP+EsiCf5G/8GRHoywC+JTeWft7Pie8kghhWewqKx1eBPYoF+
7IsASpilBmFvAOuLRXODULcrYIYQugWJSxVNBCKkUz1Mhm7cVJDrm7P4YYQhuqLtW9EDOHQBXVs1
DG2A4hjDr0XNsBqYbvfSwTPTOrZBNW3lNeYyc/PUduaGs/VfWrgjnZ6cvMOef78V6yNZjV6aA73Z
9yKO9HWgDoAhgo4PDJlyLIr+L/aLgyPxcsH8RR7s4ma/a76RqInrJADsRrEhba7naTMAXX6AXMmS
cNFddcAy9CAlJHAbyqIOJQWbyujPP1X3ev3Mf1+jbtc3kZ2I4a/ccS1u6Q2o/PhTxEbSZbQWPt4+
ZnGhtXukI29V1zIb9yVb2dNyfOBwSkfP2ShoLogs/8cbwwvMQF4OFK2FIv3PmySrb0Vho3+Zntbc
HsmzFbrZYXaGrfj08Ib7IR2bhrTCsp8iEJFZmpdFV9RzqkU3vGWj6fKtbMvzU+j1MzEPYMq9lb2x
wyaaYUWlVZ/39wKzrkM5ZR9sWkrI9BZKyBYSH8Fp4kCDJWhkguNWwbD72mrD18vh5GyqYZPV/iBB
IskbBgJZpk0heal1jHsdj+9GTsb33ntfn1iqSdjGhlzABH3ikp+4DAiqcQS7YtRZuISzWvtJNg6a
A/q5L/Uy/wL/QCKgPfk/HdHPrD5dRO86oZv5ta76veYUuvcm/ESc/NJkkblZm7qpMGbpY8Nvsr9c
AWQsmbPCsI72tBdWdw+MQQoQhzqdXhWbxfA2PXD7o/rGopuWavJiUmlbRUyggJ4xVgnPcvhee6qV
/05dMSWgqGxqoV+RBtUqrlpRPGSUJpkkjvUs+0YjdT6Bew6P5Sa+gffReupIZ9o5d7cKCnRjdsrQ
H/JhfHCNL7YBahkWeUSERmLC8wykMZfW5Oen/p31Ik0hg1ts3u24hv4O/cAZwvN+BlD7h9FmdYg5
nf97Ur2eFM23xzfnQ2eVuJi6ja1UujlrMxR/0b4DbBQx+yXwcI6WgTMwByboDNX4q6/WMCg1NHII
SecQX0nWmFLURpBR7AQMofU5/9ZZYwDJVt19iC6IRrRhJ87ggTgXl2T8jXF8h1L4pNCuQnXWQMuq
rMXdYmkNlkPwyQAJB3XWqYwq05kBEZfEXD633cboOGDS9ZfxxuMfFJDCCNaEHH+zHzNG/69Z5hwq
PXZXbMBV5B6HPKJHWH9muxX7DTj6I4k5Buojg0wylQ3bFq4YpOmefQtRFdvCgaJirsbyfegWL8DC
5yI9MfqlNKVPS+enP0N76PC86cPTYYyAwbPgtF4fTHGM8Zld/oZ/tE3wNAyhCH2kgNChgL4hLHgl
O2PXZ8p6K5/nDMD2tbG8oenqnPvLM+QBUmh1RU+f0oiSd0ott9dUVqzMT+o3H1ECksQIVkGYhvSV
GoPAq73FzxLgKxhmI8VAaY30UNWINTMSrRRpx/aPw7WBYzZn+VXxFvomxrNuzImKjDWG5u/Dtu2v
4P4MQQ4+chQhtsZLysbknad0p67B+NPLXxgQz6Ncete124Sd9TNKDQRzuWHFfxANxCX4aE51BJjA
IRmF22Xs0L6jI5Q4hk5L8ePGLp6aMfSaOmZSLBg8UOXhEqVvF/nSBEbvIKl+GgF1KWOHQvkP3+Z8
2T5RFgyK3Bnrb9OnxaooUT5HWHbQSuczH2ShhiSk18CdajxPReTbPLGNKKQpb0+Zg7XM5V10ryrp
cCnAAa7tv0/GfW0C1ZD4hAQlAzjTDGDcKZE5uKUZ0DP/9n+QjesyO4odZS+/Uxt11x95ZrzGCuwp
lhGY9yC/Acwgi8OU2kGrz/qixFBq4k+F4w8LnFB9t5ch2DsZ/y2rpa19/7oQDky5x2X3iN9l261P
Wc0BZUR6EkETPI+AoG7bWgFQwNSwCjBrKkEhLcxnXKgJ0qIR1aHw8FZ1UVckWYNG8njXXALJjd1Y
ZtMoDHs/ckAzRxHeDMN4bxS6AyZ2QWa9MS77FIO1Oub26hsjmAhcsDRG/RT1E9ID3lvz+LKjOo22
1Kaht4N+g1p6LoEw6VEkJc9tYXfMQcSYL+tQMAornYKAKZDgznNBmqYsCrnYDaaOfbkkyiWzamiA
MLisSZx5K86OpcQj1BtDFM0XOh6rMvuCrSEwcDXJMkQfnZaOJYIqyWjN097YZep+rDtscXWYt6N0
rkzPA3YjFb4SKr/jUHqu7k9Bmt48f4L4AKImvxrs9baUMguuAdg9Z3rIT0qU9py3GP2EN36ET5OF
v4kywxu/ilMjtOTc3bhmzQtC2zop/U4+2Z0L/DoElS5WXjoCm33fJGtlInsfDRL3pCzwsbr2d7hR
0T3JnpDmmj5a6tTwOBsU0FcVrz7waduxNT9TNLyK/oFJn8BzV3a9HHgJOMD8oD+6wv/cpAENfuXm
WNwZE6UNK7uZSBR8W40iD5kIg6+SKmAaGA8EWn3tATmLT0w6G+v6ylc99XCktFKRDWErSBiNzjE7
KZlz+ghaAdHPb0qPjZhlXrWjhRS0ENrkfD34lytwu0+LuhlRI9UcN0UeQzbPb0jzKbpJcMOoiCXc
LE8Cge9czpRBY1OloNsnnut8AW80uvvg6TOBiNjW4VVg4+PjebvexEjLdzlv8CqPB7EU9RobXTV1
cIgczXWDoarLx8RCcL3v7mAZ0lRosncrWPw2Jx+gSAFQyMJ+IXqpE+LKzYH7GUESE1Xszkcoxv+v
nCE+ZijlqRDy59MUgQ+iH+5AyXmjbi7c3nKBYIAF6pWSAdg9ZKe1fndbdA0K4PPxsWIL+1CGzc9m
mu/fCoI4CTSqWu4kJDdAYbOvQxQ7cO42Eh14Ui3u1yrhEReY6j6k/o+JX7JUWiXjHhQ6PGS8bGWW
kH7ixi8CgOiVfPpg8Fbhpv0K9+AEHZhCJ6ewTJvmh5IQrUWmG24+i943ID6c5pc4UcHJuxG4MTcU
LV60D5WYIsN96gQR2JfMvU5uh8SlNuHrikGYi6of3P+/BGnfEEGwLV/0kfIwvVH6hg/fwemK7vCk
iIcSRABz0mM635vzTGMUTsz/mjb5L4G2ZRog1lsRWKOVFz4q98GN9axbxkEGmXjgYmdFkv9AOfTN
JYh9Fr9Ol6pjxmOOT23SqYGoXKsY0jYwnqXc+WjColPPEwxGGNcj0YKq2kkdriGZsiGQ5TXskvXr
qfpQ7WQIEF4x9abzG2CFKIfLqWdrNzJvI0wgstnniIOZHP+JOxp9NoRCDel+eU2L9yYv3eqzY/MR
zuT6vRbTkjDwMB5CqLpfYiD5IC5o4MR8sta88HJ/G4fKSDV2uG4/RX8aPIVnsWAByKxqYB/FGsJ2
agnh4QDAMtPcUlm5Nej2RJlNsYL3DjXbV2P6+rT+ecASQJx3bUhAj8LCcZJOmcs2PQJlwnntdcTZ
yi1pQB7CIegfB46l34dimUDCBCfIWSRBvCYfDkO3Dsv+Bijm4dxdPSiDYJa4sDB+FpDpzM3qXeBj
k2WhDo1Lvi8p+8F5I2eULtF3/qFPPwIIyazT4POCkGxBU/+lcWm8GjDGwX+26qF1KyzyuUtt4Kiq
vvSnc6R47pRdgXzultBEypNM1oRTmboKLoUe0pRpcKxzhjdZ2b/fngqNbDJXkPWEWDp0g/DVuyWL
ZNf/HJwvaYrCKLxxjy1xL2FZkLF8K6S7cuF7/4p8Kq5dBD1Bwv5Q55KHT9K7TE1ymgTHdS8NgIXu
ixH+FofBaiuXXsMdjlbAs/L289bwWix+kdKo7U0Ct+FuU3MhMIWBXEMwsCyysfNi8GYEweU868jm
9VbjRsjn5Qv7ok5uN5bTm9hIF6UUsssPhw8v8m7iMsWDLPGXZ+h2LgARFS7P7nFFSEovOVYAAJxM
tmxDm8w/aJeOTTYBahDJNrvgQL8KpwN+yFHAoA284FK0G7B3YNIIBwnt3h2psBT9IyAfFamo916F
6l7/s4QOb/swuSG5kNOSh+rYBaz61QMdWffdLk4aKgb+4on77va3ggLkj+2KX6K4nSz5EcbSHEN2
x4txgM05ySamd1qCeX7+cqGbKnDvT6vyFwoB7VSw6P29VOJlMcmjRvY+diPUBdMkqiIj5k2dmdFV
5Hs5E/c/S95Cstt5D3r5/wLl2YYip2BJm9Z5FpRRta5PVuiCcP5rcyjN5rJqyTCkm/7SCg8SfCOs
o3rlBfR1OWTDxi+aSOFlh5yFD+84Ad2SWk13UpLPlnxy+MHAcL9XXYu2+jg5PfYzLfJtNOh2Gg5o
jNnE+7LJ/A0B54eHZ7tYZgwGATTy5UMiwBdfyI1j5Th7zGV+GGuI/5T7MEel5tXPAfAf3FHK5QiT
alEm/00BS9Zy7r6HbiTtYuWww++F0gtXjKPyUxScTIxOgeGTb+k+ydkyE94xAxPBJmDL4FISJUvI
fjPyKYrpBn7reG+qw9DPNah3ibUH4kjKAFMJr8NqXgvBjLeXYSudJsrdzo/oCpm00iQ6wO8mre+X
98W2zHx84GDLmWRufmwZr64KlGCfJ4WlqJ99CY52bQzdpijXVpkhoNzJNOJD1FRkvv1EUjyA3Cqt
s0wYRUbAJ1ImYLUR6c6jZcB5WCAmu3ZK1pSurWVMqESHYV9wI9S4MXh8/kZ1xL0qimRAdt3KnUht
cGuXjDnS3YBeieiwh88ffm8d1jYKn7v2Z5+uEGCsGbmDZEj7vWqadIlVk9kg5L4ObW+Qc8zNyltY
xfPbyCQLTLqB8es3XZZb1i4SzW5OS6pcMt2TPg58bkoc/d+qmyjm3jt08XCdhdiwSO7Qe5ix4Gja
pO142sbulGYLIWTkvLUo+r9QSmZm7b2ncYeln6jbER0ddlM687rgtEu8VBCcYa7KD3yFH7heHnsC
et0MPokVMIAGBWJxeNxAG/cIyvnk+gk6Z+RmAeKq3xSSbDFlYBXWIK/gZ6KjB9U7VzwFmxqrv241
dAbpXcfK8901kDXxKUq0kZ3BeRE/kpiyRcc739Xd7JRAgjzORyWmWJSxTZmmNpyiPQ68gZbUkAn1
xvmrCZYVDZWiWG/mt2PiLM/SsKbdcwCwX46PUcNUcwb57TZrcOelKHDlmU6YyrtCSPG2oTsXut61
HkrYsLdDVlHUcVbPyfiMKao7ADc51BWPVx0OK1YgN6ox7peOvgpDUJM5zzjX+XKzHxziVIEtBQTj
UZ3KzMXBtYJjnoeJK+wfteyGmPszLIGUHaHAJr1o9IF3dlKnbSdafvpCjqCsZxJ5FHlLfzP8n6eJ
rPVZR0KxL/E6zaSu1qFfboDbhZbd551HFhtBNyPtBzuWhGj5yYv1ghtZUdYk/yqvhc7EXAeLFfTk
0Lg0WdDysKHWaWeoJPhQUZkbzKJ7QAi6C4TpmVQ1egkFIPmTtXU/ZdDFlj4DC66FoE1nYSV9ByPB
AeYDylUISubWukbs5kts7ezM8Y0McG5Zrq0dEowPew6SZ2oTTugOcwfXwSX3nITSfnBEXBEhFmr8
RusSejzTnak+e4A+BLGmhMdNANAs8x9NDXm7LjfA9DLu38Ae+ei+SdgYCVdoDydEpDi/epB7WPk+
grurlHCLT13A65RERk9Fbh7A6/2w6LYBRyQ7GZ6MoDx5oFyU4g9OhsWsDCUtw+0BygYQWw09KoCc
3Fql2isxNBc15fw5MC7LWylXDgoKPiJn/kF2BPJOQWHAIPqVxLqJaTUg1R9nIhZi2ZXxGK61Pipq
IxwksprrtAXA5RdVJMO8i3rKScCgP/npBRv3Bdv8PYCpCCrVmXCs24mHJ+safL/K9Ejz31QiFKUT
adTQGid5VGQl1SsRlHyqHCx8meG3MM+N1gyBCY6/RlBmaQ6QPXfHEXDfocVpnau88qN+L2E1aGHx
h/0uPfBReWxXH7kQeNhmoxbCdadTapv6YC0blt1wXxB7TXLDGbpfbkTmyfZhB/VqVSFsr/OpszLn
XL5Fqn56jDPPADHF1G8cN2xEyAOOpwVWFYJEyiphP++qlVR1DDlFmglCPuOPKFmiCaZp2TNsmRKl
/Xg05LOIcW43agLphskO/Cq6ntQ8J83yKwqqg4L7NDfp8mLJ0ypFXQfQN0iWB1cCwB/jCmZL8lPH
EUAos0shcMvgygSCYP/5rvMYdfdJpn7MbiK//vgtEf9FEe9VOmTWAcN+AE7OyVvIZHK7iqKcJM3n
LGAsCpGm/jzC4z400MoJ1eEXm3VRTCncSORpXwJcgaq7WCJ4dQLOzZ47miX6qPIilpRwidu9t+Nx
hDX437xe6XX7ZOYyTXLwOyS0HU+0jj6RRIaQRKl3TGDlE3Bg1rn59jFdtL5fgSAe8vYJ5GMsWuHR
n1vLOuCM5Xi9VLQJrj1uPgwkCzrHz5TOa+LJ9Je+KXEMZWOvZ66QvOLKgs6kXQPwA+e3AojY1mYc
jUNvmFMWNNkIBKPxEAU/W8xh92iSWcNNFNNzGAjS8JFg8EFUBrmqGiN7C75nmPrbqR6Wz/EiNQoT
/2OvQYwUBDp3WQuhI+GbJz9i9KgToKhYyOwmnIXFvIoFVpP3kRBPM8l7m/IvhdR1agxLcA57kbRn
XMz7K5d2iMtg9Shf/QnEWeNxbdNgRsAdpDUsGsj/NFKcSfsQNGbGGlFLcduJwfDbWDvDunMUXsDl
xEecgjMXefUWNVq16iRDaKLmOOWM39exdcR6nh8nf60ne924hUdtT4/vsUeMkK74Mt50t5/8p1xj
XWn4SA44EukXw4dJvgwFdbdinJOAPRuIv7auj1OzUs/ndjtXQRupddrgIDp8gihq3WdcHBPgxmrv
/xCepRKmZdVIngllM/kxpN/0SQWsvgx375aYvPQRRQWDDPAaRKWx+1c+FA5IrrT80jwtbN4DLvC6
JVIO0sMvP+x1scZR03ju4VOq84ZKmsiU0ThUyNmgPr0iZZAvSmbK543CKZFNlLotxENreH5bEs+X
F7TYRsWdEY0qWcqp5cLb7psTnbHA6Xgu84gmdhimsy6KXoXkkpSVEsyMu+gMLxCpfzA/LIER4iSU
E/GX9dESeyXBM/P3txxcA7Dv53yQEkYmaP/w41kOWiTYTdj0uXznUHaQCnXQXfbl5+ECy5/0OUOS
eEZf1bTR06rXoYQY0pB7TchN7ngTAppGiNtNZPhOz5oYSp1eq1t4gab1fWjlaZkKDFFpmPmR8Kq7
6ev0vF86vR9FtIzRpWaKnEYfxhQivzedw6wJ6+RgjaV+dyi7beLov+UpWhFyrecDcJ7neFqjj0A4
RLuBguNanCD9wivQTnxB44nNNDNSt0Uc3XzhHSXSlfz79kLIJUN6LurR2k7B37KwkXvyIbgO+2v2
rlFsFH1ldKMrsQJXGE9g4950Jhe3OTm39L4zdQlHGy/8+x/OqRZK4UvbNxA6cQGemYLUI3JJFTjZ
I2CYWXNDjvCeyT6KLsgLxn2tCeYhyzCuYqKcYVcWq8N7e1p4F+et8KLH0boiFy1qk/PXJS9aITGF
qLOTuIM+j+3z4Hjyf03tIlv7euwW4VWOcsiIpv5wCIGeN8HdzO9Qo47by2LpKo8Z96ZMfDK+Fcg6
Ybqn29nHjrsH4E1iaSjzJLUbZdx3Vg7e8DRScaXlPi/1DhX24/FWncMDeBYA27alUAN0SBIu/peU
dYVkaj1FGxudAD01AXS0eNL6GesDt+fuhECnCdhq9cUEG+Ly6PGmdP4DDPKA+Tnd1yTzf4q8300p
3DLq03Rz2NeTYy5iIUUXu9uqH32FC3gz2Tr+9aFq13XsbKdNZ546mJYJpdFg7AysMlSUSUZEEnAL
fwrkhi8rtkAvv+stgn5wnipBe/lmY+PpAqDNg0cvPzdQRdbN5ZmVqxh7/xD2yrJfUtLEHYA4lSNy
VWXmd073BEjBuzbZNGchuG0uVvcZFrCkrQ+mLkENC1tMvht/5VgNcM5S9/o8bzTmXO4i+BhQ+tbK
vX3A23Ayr3Dxym8PEfoatkhkjAHUA6pexfLJAgpb+EjiZgE1LeLTOFsrHXLLjqkkSpVjShyo7EOx
oRmQUrW41LJJ1Ww116n4nkCloElIXLf3dAJ2yzn56jFQcfCOK6R+WZP62c/EzxgaWUNHEM/yTWd3
ObKhv5Rs8bXHBmGTbgoMyqcU9J9CKeVfVU9IBCczeaRKQ3m8crn7NVDaBrR2MBesgUCWO322vFH8
wPbmPsiYVwjYP9M+k8GXcKkQLnJAOFZQ4Wy3X5pC3vwo+UCo/Bfn7iBinETWMq+CmtzTJHj1rrnf
NmKvOzEG5CJd2ImpAXToWxIFDgMKyEah9bdFZmt4o5zqhNL9zDzfhZdek7fFAuCtuBjGQp74Wk8+
WG61r/lcflUr45ugXm1cuFdabS1/U8gsg0U0Bvzh7Z2gBsI+O/e2sgtFqwaIrNZRCK5CaDXSCkVy
ztHM22vvTLaPc+kUzqpewgMewAU2S69K8++p3JAW8FGpmb0mqP66IZoXAuddCk+NRfKpgnkAZkHg
87DSq0qm0sgYmzXYEJLXGyOiU9871S2SRGINSq/zJSm8mXSS6iDRI1wwznMT+PCO4Twxy0/Efgpm
cP+6Mtoe4wKZO8T+xZF8301k3Znsy9wVkh9b9tsanc3rn7so1shq0OJGbxpzTz9II10UOu2+bM88
eeoNLHphgAza8iPALZX7AphK1VZbfa8/XZdoLUVheuoAt+x66ncJh8S2x9N7BAujbPZYkI5boAz+
QCMQSp2R1KVDSa2CfqqHnYjRQLdFCgnPUReQk4Zhq9IqwA8ItTv3pqjo1y1jTLstMIt48oqy9Sxz
ZFL5MNmbCZ1NghIdfw/cUG/Tc67yq4t4V9vdb74+gb20a0Cy0jC9RWJ3lgcD4dxSugur2troTNij
5BSUecAqUg1Q9lZoxN5UOQYg5F5aKfGxFcjJmzxxSPqx8nPeOPdP2Pns04ylWfyHg4zHMy9zsM5g
zRXEgo9UJOOgy2gwYM/cLxsCBt3FMC0lPuSEzdXBxh+4JhQHa5MJFXHgVp7SiXVNEnE6UNz6uGSh
9LRfg5EWOMqYyScC0W/3C9KDfUSYMfh3BzZ/jQmczFy+lnAHnf2e+gQCz+cAFFRWHgTKkVlwT+ON
rJZOSuA4nnOYNp4kY1MVeKl6eZazibkEbYBXHZkaLSVOOpfhR7Ld5AxJ8zL7m3aVywBJMYQ/lin2
byM87Q+m75PslrV376Kh8McsP3Ai2y5Bc/Q5P9Vf63HBqh/b6+yBoa/wlLu+yM8+6Jytd8LsWKaD
0eD5aSO6xONTUBvKahH0Zy3IQFtEx+1vzsvz7IsZc0/BUx8EBUtGx1fdE9nRMqZ/fYMX+FPRSrRU
46yopB+fOLOX0/AXrHVbpN1i+KvQhccCRaBpHDdtYz12564YcoPxH7RlkSf/yI1ZD6r4oUL6dPeN
CfZhW3eZEP9RMytB1px4GP5Ypuiz6+MKi5qmS1mB3nJbB15JvInMx2ktpCjkw6uBfJ2aETOE5Dtp
eXRMqubRBBP/T3eQsWTDbnExf+j1JR4vjXakAj041PP7rYRp+TXlKuLJ/p0lyzoHgVaWMwa5eBtS
r/+N4nxNU4EcM1eWTo9tqpUKncPIPeMoxddfiKdRFhqcLNxd9IuH6nROWzWLNwdVqOI/A5u3botG
bT0iRb0oGwUIRONimm9pe/FVstFE6w9hUDnqqwvX5veIOISnE6VXcluxfINlfGDUOJHVIrt0pMG7
nepKfVpHswJ2TR79ruoduPW0zFTH4cVpSGRqDvcbuNCgzHGlF/Eg79kAE4kBtbT4riTslCXuny3B
BJCy79ofUfvXEQnVjEHwLi520xesYo/hcpL45d/wuK8MLxBbWBC1IcsAe7Y8G4nEeZdYgg7gj939
8WYGNL0UGSNZUaH4XlGHoxoF4ZiDEZYwaA5l7PHjaJBaZcyan5NJKKKZumyd/W1HzNFGeLE/uxEN
ItRURrSWOB1h0O5F0qGaEIPNBPowSHMx2c0cq4iK7r9J5PLf0Bjpnh+dQmDndrjTWf+JRXFHTf5H
b51HnrXA63+IDMxflNz9IbJnZLYxjzVHxhZt6BZT1XxZf9NUpETabLDOZ4k0Q95sUvGdO3DmH8DV
zzTPzUlOzZo5t5xV8VxcSvFta7eairtQDDdQgnynwP/Of6j1W68O05ME+Ohin/BUnlriiJ9tVnxI
G0yB1Fuccxw9CpKuDHZNX4qpJV9PkfyNCOzulYv6XFlPyZAVW8Q3bzcDnuhCgDbMwmncCjljb4XX
sq1jjQVB3ZMWFPg9LjT0VlGaOOu+pIy0z9mZj5MVyQESiAsYtFH2d+WkAg+n5+RL+bTwpzRjJoxr
BWuaaYn1GaMc0HOO/r/gMYk/sX8N1SWEim3TFIuMNGk4tptKpjzQCh00KTQmjQa5E8bMqNUllj+B
ibRk/TLPKnrMVC1ETxDTUGl3zDxvpOkW+7gNErst6jWuH9z8mOtc7FAjPb6caYCZdcRE/5gXq2Hv
lGLiHnL1UQzFqqdniS11oSPA3bMsJRUGUfgecU8kylsDwjjyWQl/izSGptl+psp/5u9dhHhf6//y
YZaxYH+i3Zam8T1BgZVLm0+qsrjwoemxrckJltbXCCXekvvWuvYTfT0eIq4kMxPOXX6acGIfeiDl
8rv1siZFv+iaGTdkqOsAWqsueW/ww3kk6lF65jgHahjdszgxv0AjZcFQU1dK+WM7+Z9p8DveiTQk
XkC53Z5n60LeOSOIL/PO5O9SFTMJxE3AgyYR20tXLo4i4DK6JvcNXiCBvI4e7a4qcGh4ieZFZAi4
HKnwVDBo7K/dfAULvl6GvPcw/xcff/RDZDv2LMIhMBwYDy+YH8yW2HBvG38gch+UgYr5wBP7zRXi
9/Hv0BQyykgdk7JHTCRcdvyqA9ZCgDatX0cRFAdFkX31zkGVwomjDFHPWS1LImEYitfHiAdtkM1P
9WAHL/nXnYgJ8huKnBHzZDw8ERvd6qZtFaykgLxvTQMtEMQuFrqpXyzmCxvi2kqP+Z50ZXMeZv01
3LZI7IMBkkBl77Np2dxchCWt8wBDnCBc1EhEexIJE3TMrjoInYTyHrR34KJWndU1u11ou0wWOlbr
lTFNLZIpvXtp24qNzsPO8EuO0JR99XoEerhO9prr5l6DkPd9h1wDf8tlgmnIlO0cEB9qNw9Af8FD
xue+AUvwZ2VqRDl3kwQ0off//yCgHlVOXUYT+VQir+m5iKiY2oNbNXn1T8/8rJxKGFdodrVfWdTX
nUa8HH7qJytV7xxiHXN4zTS1MxUrVBz5QY7/3agV6bQxsFwsrbjwZE2nQlvJUWdtaq4dUCAC91o6
GDM1rUHMaii3AN8A/j7N1023rZU05ZWLK2dCdLahTWgku1wBEnXjqmwdePUPCEbbumfo+A8TaGqj
gjRfkRI2gTWutNfm0C53lgAVgORiR2ZwJx43gaChl9d8M9qbw4qk7QkgWURZDAsukjZ0cXkm0uE6
oZ9rLsUTg6/eT7WdR2QNO+H6zyMAdr8eOOntB2NyMEANJ9lwGHv68XSjGjwNNauA/UN+ImBGCxvu
jUw67jVTh4fPrJfUsDJGRfkesP1M0U9T4tHenrBGAa1Q3+v9PZJj9kum/h3Uyrguj0X01aSy2lx6
d5a/Kqb4oQpE5a5WkWn4pi9XeDRK9NmBuRAJWkduHs5rFtLqFqj4KjQOqDWPia6Y3MkDZ8XadMft
WGIf/7w1JmlOwve58nXomsLVSUyAF8IgMVXZ3CH06EWTNytVw1qfd9DTWekdtkl04JbPBHNXWzFv
ZbFWHbsWb3oeWQtUg7avRYdSSr1IMNj7GUzwIm/AWVoUgHIpR21Ns0lR/xEENiTlTnJ8Eb7cBN4A
E1ClTcNxzPMKMiXWIiVtekum7Ypm7dUvoX5aZ3KHyYHniDtXJDO2gLQUvsujN5pM4HZh1hk4HKpE
V7drICF85WUT/eoMI7aOWg2M/ccvC9VXK97mXfwTollE+YLPDDOriH818aiZ13xsXAoZYKMK9gci
yNv/1DtHnS83iZ2r/QDE10/ANUSviofL+lttDCCpfoxmn2WAvHdGPpwnguK0tmYhBIsAmvX1QXMJ
SsbzT1G/mnyh2me9seTRN1EBaX6plqiiwBJy98alha8hqr0lzTexlvoujVoodYsbNX+IHQhUnMX5
RoJM2qQzshc8R2ivLlC0C2f9VC0vfsIx6WaB9Ci7KQcPOydy54xmHUd9oRX83KoIazkLRonGGSXw
SbpvBoPd2GHxwlQZ8n0v5ikarhionf2Q5KvvMRcyAlEoE+NlOH5pdoVbslQPqvnTabnYJUQ9sceP
iPOD7stgweG6JM8bGMNTHPvGdVc2eC/UJYH+YE/SMfNDP5QENCGlXn8JGFC9S7/qFO1L/uZ7LcnM
NGA2hEHRyNL/gkgyk48sj8UflHVnq+49H8zqHp+EvZP0HF4VGqXNlpVtPt4SZDhg/KwUWzRqYd+O
xID60JPjoLvovbNBD5IvKpMZeTM8xVR+gLyNoeIJVM+8z7T0TtWFKKRjnywbQEQu7SzEfLWU3L8i
2YMX9pUAQH35IJUvFTSta2hpZNIyw8tUVWBVPaWK9DS/eSqxHwdQDnkZEvjSfOknyF6jtvuMHc5c
w7q+B+PDR7MLbDQynu8aCySoJYoAgI4yTN3of5lo0pAJMdzzHEUYYpV17S9tKR7YWAj8NK2GiLf4
Vhq0UWxuiaGFazZyDndV0uLwCzxm8HbhkeIYnwp1r5jL5fwPd/FXvO6jfP04yDEbfVl/VZUViHsI
1HN03WjQIzTjn9FJrqNQssHrBQMNxrlpvqCw/ZjEpCcvMcKKlJdZwzCXz887p7c+scLCZGHoar/g
IOkEag+eRmK12eZMzE5XXKaIJ+1vLrN2yMB+WT22L3xlCOs4AIgaLXhE/suAByAwWQeBKF4YU/+k
B/5+wOR9GzuNrB4YCmIDrdEsaTm9oYr8NpHlgijphlttzsAOkau4ub7rDVA/J73n+ZAUCyuzXrPF
9TUNiqjMFn1s3Aq7ojHPDo57/ACjy1mnC7+djr7kfCNq5YYtnqRCLqlvk++SE5bWT1EvMQd4KdaB
U5EvhJTlNAm7wuGFz058F1nl8ASSJFwq/9peU6tP6SLGoZJ/xvA5viUygUAjBWHrfLhtyn7FrBCO
2ISm6GWvCHj6fkOip2tmTUReTzLfrWoniFiBxFf8K0ZJEEwnM0q4hOcf1ecjNax1FxJ6X7ALUCBh
j69kTGBSlKO7lLpFRAFMskSs5t9VQQXn0kc8vZUBfmq2X/os4NqTBp8K0MFEl91X+bU/5Yg96nyw
89obyRDnlVLry2a7eGDGCmnPsohsKPYoo92oep/RNJMyY5J/J4BTUDX6teXGgMoCYcNI63k/0b26
0jnd15rbdbI9UR0EJJAkLsdmlnMfKbYLKZcgA2/cXZR7po4UmuEvHCCpw7iLy+RSYO38euh083Y2
tWud6X8vbnwZBh/7ZZ+47i7SzDmjFCbG+IltJnj8NPLEIOY/MDE+hRwWorYo6Rv5C63pIFm4Mi6r
KJLyX51+0O0SY2nzm1KvIPZx1UDF6USGh6Xm+q1a7MBuHdeHbzp6kWHWbLviUeXFOjxFbnTZ/mEw
zuRjUVhglFVJnWD0ssRwN8+J84MXn4Qg+GXAwc4fVBYTWGtufX7eyfDNvr+Ah8lNgrX7S8L59f9u
j2U/ccLD+R6LoeLPWSBPRAsj9Sgm026T8hYx3AaNQbrhCHUPZArumRWl7SqZ/4oKEKflp3+eXCZI
cOC5G1/AiZOBVxUY4FVpRseVFzyaHCg1W+HWmwyu+dssSZiHKARYT7gCjK1eGjJ+EvEaKh7ajUvJ
AU9yXkH6ihwNVEO8wbNRFRAf9coaPo4G1rticQ5T2/nso//GDDkSj0rf8OpcvzIjm+LGiLKq1cgy
DzYguUwE8SmZrn4tfqWWAuNHqlmpKd+ZEa3/PGe/fEF6fA+TQTSiYB2u5/Sy0NKcTgKzxkR4KRsm
4rdLgEFpaGvhSm0tyQ6muEf65txzndiR7OTrhl+O1fBDQSqUAGc+q0Z3exqK6CaZc/AXSlYRQ5HX
BkgIVMjvUBxBkK6FleHO81A3SPRV7NCQ7tCRy4/CoAS5wtVp4EqdC+yEqtLMsObFhHSiSSanFpcN
99SEX7ny2KhOa3yaAqGTs7boC+gmqh04W3dqL2oHrjIkqutZBNn/PsXtBUxzJ+AVoQZbEuuvl2nX
/j02lEcLvxKC0IVI30Of/CQ5EM2bksrmpcwnbwAh9EKYxFMsrOn7mhC5t5rfWZDIEk6O1RlKgkMy
pbJhesNLM+M7ve0BREi7hzhPY3hNwbc5laAvIIJxw1dzE2nP9Dvz3BqcDC+oQoNdizomjd9PjKpI
0vjLH7xTKsb1qfgjdGpl3Flydc7ShE+gDuadin92/OOQhP6wfI1bS6L6w+iAWCuAeEk87drEBmFN
YgmTk01Xokm+VD98ZNMz/bWlWRqFySdNRmsHApD3ZyL0f2QpyKwVOAUEMo9vVtepF6NP8+4paQyx
RSwY3XyaHdOHE8Z/e4yCS+Wzif7rE4xufaqRUYpjJzZGrWA8me2XelEwSYS7yK9k6GjaTNr3sDff
qqOovsvu/EPEOULKL/LlJXE5kWNJ50+RFlDHQLRN3MxwSCSgEMUtw3FcKmeDirV8JAASlyvr/uYY
wTnmqQ9BKJTE6XTLdTE7Iq4lhOD0JFXezhfyzPX12DO6YvAfHmrOpcSFmI4Z1a9D3Dev3fx2Tig+
ps49Y6dCtrtSSd+RXwG9DgIzUhqRp6cuPTqsAVp2zwPCpIHuu75i2nFdfV/XiMzgCOODcEgqHPet
01eaIsk1solElU0VGTJ4pqjanXnFTznzfkbGL+rDItBEfw58UOIn9j8LcmVPL9lHoGtdC3g5xlrx
0cionyICkWbU05XisGbcrlLpsSFRO9aFvK8b98Ntjh+r39qvyXcLTmriQHNJNl4n/ZNWEXvqHACs
JGC/1YQql3MCCv/pjwK95u/eP7Ggw2OC0mBjBj500AQVm0gaH9gl8+yqUCZ8Ijr05zazyXzp1elI
NIS8Dhyx6hG9Ci1GpHSfAbigpoT9kH9pq4mwsCWa0WhXrNlc7Dv+yWsb00rupsHWHct5zCPfGAQV
NNyjTENH9knLkvaDvGCetsucJn+0GFTFX6cmzPqbbU4TKWhO7rb102VOm3VAq65vKLa5IYomy21K
i0zNjBUPVbOgyEBC/G6/nHqflXbyL8ANbFvcPwHzmjGL/t9TTvQRB0r+dgIIuIszD4/BMc5BARbi
65QKlLegioA9MTxmWaSeXrNayYFCACa60SUbMCDFokPHMy+stC9U3Zo5Hom4NPeLDYM5Ng1oBBff
4DOf6xxDtYIQBuGK7zGK0e/rnuiVvVBg3EyoL0B9DR0RT4L9yehbdYSJ7+UKuzjaenDy9RVzUJrH
tCmOM0mx+pQIiIKDJzKlQNZ3v1qeGzCmHPQbccqZF69LHZ9cWA+baHEEQwtwujtQ+Ur079WN8FZv
tAZJcHXYtidUSd4pqQGjvJSueJ9Gtd+62KrByQmFV/xI35bToS170k5rRa50rYQxAwT4S0rm+u0m
hzMy1wUDkZxJulJgfQz74SWa+YvW2nNP0RtH3rR0DWC1S/3IYKHYA0esh+BZjwa3TXK5393alO6c
Dj3TK/zs+7XmvJEIUhrZBcSVex96W5R4gNscPqxmh+D4HpcwuR9EUeHguZWGrwavg/3ZLsqPjUik
/IkB443hzRJ6VVQjtp0GR2OpMc3vgdhbhQALUKR/TlUMJwk76BgOA8uE8u8viPLvijDSIF0Un/Td
D9hf4fNd/TUQMfX7BKt+RELlcgP9wy7ppnPmyjA5tk2lBu84hWKE1B7/Z+u8IWNewSm+oxTpLTkW
dCIVqWh4vYmNYH79mwlV9zmf1UFCOq1UBfydRWaX/aAlbM8rLTBpxkopBT7VsNH/g/a1r9Mdg2lT
+arDt825qXHtLyVrJxAgaJiDE/om3zVfM162E/M5XhtUi9oiFWfnRx9WSfP7JA2H8Ju1IXTd7BcL
7ikhRK4UOJTc2CoJZCIV874nFWWWrHeKAIMYqgCU6exIuZGypj1dUU2mtcvCL4AWNRz3QH6rsjR6
/KsA2gwig20pUTy9qGWeI+RBgyM+sTmCMOz1kqkgGuKCUa6kmlj2uHeWJa58PDmjKRwFrXaVbbXg
abDa5tIjTrDEDOivj3kzlIjIuUbGCAC2H8hg7lVtjtA+gJ2CDcPpNQHUoSBy5YIoK3zmgPEu1NTW
KZuAtYgLdTWvs/vwgQh90kl1bZlmQl2TeaJ2g+ajMMbg+tbrpEW2gxWD9/BE2JWFNfA+UlOc8QSc
qhNLtlzBQK4MIQ3tRiRhpxYR21u75ihBn1yk33qVgH43GEm7Nc7/TLK1m3LRQjumv/GwtWZj3hlk
J40mNIwnbRUVf0D+N5JZjnErd6ibYnchfwDLuFuCojz3E65z2Copzxyv9Cj8eA360mORjgxYlUzY
lROnyAhup/a2RnaTCrf1RVLQ/LorIXUyLjicwIknFq1IPK5KrpKk5bc2mLGUS2Y13+Jk/uVOGBqA
hilOMjT3iCwA4r7HcmG5BCpCIWKsgx6xBunSRcIVLNttbeBwCC33RgQetP8RNhywqID7xeTrZis9
Q4x9ICWcPdUG8doKb8JQ7DaykYj9QSs1C60diGwi4eYCYYGw7llbtbGXwVP4inR07MQkChKZ8Am2
+LjWXALKs7ZxoLrtobXM9I5ydEA5/OxiHED/Y3IoU2LGlgmEwXkMeHOJooXEP9kwDgUNxnpguReY
aorUqcjTClG8tOvh9/4xPxtqFBYjwCNYVLwMirBRIKNNOWuFQYNs4Cvlq1gdIuQJR7yVn4wrR1LI
OHRAcBOXjl1krXekH6mEiR3Gcp9VyYEq/yJ03C+RIo5mp216XPaj3SSRHIiVoXtCbwdj/OVdKZf3
XAAxygXoDGlPjmtuamqNEfcA0TF0+XY5Ssi+85wo5H3pXLeOCudgdwJyU0VWBigB4LbG81hnDfsq
BKli73rahyVLBqQB6wnFB5A4tNTtzRJ+lwt+p1vsqqJnQSVx35CkCu2R+lh2cl/2z31F6SpLyRG1
g51pu18Z9TOedApsjmVSsapYHBYvs90/lqyYI2LhW/eKjy52lqd5cLRpUtOgrCEdWI2xqNIWAAz8
PdZIJ+kdUDf7tw6jFvEIF5Vev5BxR1gqoh3+Ue9dKjyjgmWcv/UwP+niwK/+tUMHcvwmIwYMkrWZ
1DU7R2oCrDAw+nwldTABlHAX448pIYUegelyYOG8dPqQgbskYFIirodzd6nrGQ9LRppNcRtboE/2
EBGE4jylvJxEmHEq1/NuW1OhFwQXuysWJgXZPhabSAUXKJTbkGB4XU4DtbxFVVyRqHu8vfegVeAF
k9J5sX5enoxi9Yd2FTlgXuCc0eL9o4AB3uX77LYgGdFe6XByypzeYtMFT4VEeT7M0jovQ05HlJ9d
u4x+5OXE0rxtQxIEKanJDndokCfBt9IERRV3zjjsuA6kz6XzZymDf4rGb8VrkvfU3H1/JHWO3xSy
yV/X1Mtn0QRBGzuFpTR7aqGyjDSIttYYZ+fir490Swkufx2XRjqeri2KOeJiL7sdvhbk2ezSpcsP
6naYi/YRjfpTNi7Vk3/iydOfIyRdgf8enl/UlKvQckS18D241yFS+oPwpbxpAjPED4wWa5peB4UF
nYrnyEI8Wta4RzNiacUdJjX3k7AqFF/JumHVoeEbmKGRofzUo2mi1gFf9A6RtF3I9tvm8D+CuMJG
lYjX01rYvrq9OQImnlQKZ0P1yePfpsMC0Oht2hYBV079oXtaF2UGiHKRJ9QFwDGOvQ9bJeRwqbGw
GPHjDSEGaRqCXnmFjGSC+I3pdJKoZj9yyuJxr87rbcLHnDUCuxJ3zuAYCvqTAJnLDsgI5NedAbe+
lhAtSyidF1zqmF5n2+rFFG46OGxRXskc71M4LSufhVeFo61/YPEJScVFSAZ0i9FsQBJpXl3eiRrk
cHvuomre2PC2CDa5CJsEWG2zq2CQz86Seo0raU1yi2DxAclI1jiJ+fLySGyOzpWXizURUqTSZlRM
8o2Gb1xf2EsmfvgKQ+xFjpDLX9uF5GUJqIUWCEXOSFHa7ojXt2ZC9jucWuuCeciZmR0RBrnB/OD+
qVuMnLWnNr77CAS9EkKNMP98y/VBFSBbx3XDd407VA5p++b3usMRgMgFLOq9OyIYxUKOhaqhe2Rk
75yepvOqemdc76c3Ny5c06AMIOk+r/02jkv1dFlCEEu5ZZJspEgj2hazuE+KG+s70ubMxm9o3WgX
iAN6clf45mNs/TB3K3SSpQ8CCZPJjTEKO0mJTcNAw/Smb37kt9IIZAMfiAFzE2A8pQ0B0560rvkm
me12ruI6c04LfDeIvnMV6f+wWuCLOVA07qByDmpZXgiUuG/PMVGWvOWfhspLImReuvDEwHXHxTNe
rQ8K1OV3RYTQMC+Y2IUPnCBS2rqKUO+P8U3jRQhOYZ1Y4g0YXZR6PxHyVMbA8kOJbsvpQnGNqXUS
V2B7ejTmSILgSKSP+UeJji0iDJ5/vHNuMcoWUcBwwAy5L6ixDzrbiYwOMhaxT4S10sYqQcD6FllN
vXM5Zd76ZXyk8wwEYSKC+72LDiXy6Z1bFTEGmMcO5Uko30n0L+XKapbwa9L4IdrLsrjTFRo4Uw3i
FoZWT+WgnjWu4QNkS1VVk6hNoxiq9H8+eRrJtsiuddDa8LFDYop37BOkzRmVza6lFA37xQqOvQpo
zqtS6AgYXKh9J53FR7sh1wZ9xMIo8kIm5AcVYffrgx2tbdBz9jhNbJQyg9ib3+PZSqbdLQ/TniIl
o5aosUErs/a/B0ncPJt00NW8AV3yratkhXlJVpMZ51njEYQOJ6K6mAC4LNdQwNO5EurifPmkDb2C
1Y07D16GQU16dDgxKc1hDyBISqlhwYDguZ0FMMY91WuI986DXRh5yXNg/dO6YMbuVmfINSGLOw1z
jgxn7K/R7w0ZCVsJYXrRnAY6+pP4rYXGzv0R5IsPy6/Fl35v6y54qD96s9z2DgY8KxuFJ2fMwRXd
R2LY19hZXpOoX1SkhujN/EiwUuEZGSQ3MlZo6L6dHXvYB8CFqYUDMxy5XSsCJUr00IiERleM3h7m
4O0pftUQPej9Lp0W2NK7SA0vapaJBeUmSJ6qEHvyWGLSzzTVwyemvzDd3KWjykneIcclbp1qG22F
Zu7zRIV0jVFkwf9nnECCGTBIwf1/BCPId+oM5OY2kApRijV00XUV8UnKUMmRj3iiWTNnaKg0wz1v
8K1tsnmUPYCtkweD+ILHxwEIxPiOYXzLc839dsCNhuqfLDF9QcZnwoFtr82lxTtx4btLDyLG+ThT
1QNCv94n0Ujsrv6mxRgiTT3fFzszltki7zAFpAzj9piuXLMS0wf5d2dTTEo4GSSkIyUF1FGPIOE7
C6RybQhH9KKvxU6C5qcxOF7Xd/yiQgfFHJM8MT8GxUnRr7gG7/ZbAJ6iujzBG7kEyamMOVEJi3dH
rSidueOZRqnExkPV64vB1N5O3Ey9z3MUhbNbmWtbVdES6QfZqpp6FRDw6jzN3MdgpzIGeRacO6zD
VbXUzPEafFpc2XDukl3swQEo/dVvGuLjz52HfroIZa7bP0t3+HJPYsFhAJdj/4STxdr6vgHVBXVu
NSdlzL+NGjk5RfeXbqfbecTdGcvi1iJX2rpZ/ZcRIulpdLWRKIc3rJHkBV7K71+CxeIaDYTwIBbt
8EwJuNsvGqYtXH0h+FdvVLR4p2K65xiLMbP/Ctl50jKhv3EW/9KyZxH5VQSfTJw09YS3co+b9yip
rKivhFh+DcthHU6XexcFAJuPfLvkYHGakc4vUF5LJ/xrxr/YyEJYwNglvN+N4A8EroRfN+iTq9OX
/BYjiOpqjZy/ffqU/glG7L9vlNWW709sCWfcZ126EoTAmj5jqFo0zGw2hVCa1suEN0Jc0wYcKI0m
SJ2u7pzWlpoejjy16EzL+iq3EzWipCpnWypY7wNgS0yJvx6pD+CmC1PjDJ5Ah8VJ3w5QrPsO+VLE
wlIe6RCb4TR7IG8B8YOn/7BP/1jPVNvcHizuKhNL3Bcbm+lVD+7/Nexs8tC0SDfzYb8G1IChBYZ8
8vtabFPj1n7kVkhcz5BOOaj1AC7NFXNGn+HC6Av6E/jHiSJaTyw98o+PwHMTz77ciFjdhpTSKWw9
+qTa5KqnnPFFwP/fiYSZhai0mphIADKmbNg4e2vyujw7L1MIKc0QQRXX8skRmtT1dyiJ1gke5u5l
RXQ1gc+04bWZwHZeeF1eCK11b0ACS/7L+H2kuduHymB8ES6MU89bYGDB2PDCt7g1Fh7zNACmRogE
HHwzQZnuhi0ABF5NNi0jSv4kbK7GR6aKx4vLE+tm/SjI5ULWga3nFJb8bHeYC5wqlwo3SATNUa26
U1X0DKbqH9WRwI2r3rGfES/uuHB44ZVIlUIF61uVTkhSeE5n0BTnxFw4cjG4ZMnHfrSg2g5GLu/Z
5e5x2cJQERhZyQ6fVBO+IuLL+o04/H+OP1fURCKNmioGa3gE8FMTSerCA+SWhGAfyjI3Db4g2eFB
UKoJWtmjdTyZIQcl320hrRJ5Vn+whycrhe0UX9Ad8DpOYTPEPKUVrDKiK5YoPAs7kJ1xNQ+jck1f
UwcDJE37B58dT51bod/xqLwrrSa7Raih2ZQUhJyCZBbCvGnKvlWdHM6QmsGDDPKat4N89+WB+Jea
IJlhfYfwbziCeXDeiPUi9MA6Ph4fMcjqKtGSHIk79bum6GCgfr2C4+3znSqCTS1ThsV5pcicERao
xeXsbnvpCdF9ksjQVnNSeunU4CpsD95dxg3yMo/l0SKHICZDy+FUZ0jOMGLwASy5730hOuOq4wF6
/Qg6fgPzMFrrXb/xUjU8T2cCplCIDpp6RvOK9iJS+6L1BwfRG6x1eCyI+ljpW9I83nWeA1RSuImb
L8YZvqlWM6FT5+lNe1SSbCNCZmESmXe2S0RebNxWCA/LNBw7DvGQkyO6mg1vQY6d7HkvUCgGkqhE
NJWmEaDyrYVdVe566jYhtvhOwZbhndwjGOuFT1lrjp0beVYZXU9pRtI/X68OjU6n8ZaCIWIKDWRv
sZUQVPjClXp7iJhC7DTZdnDe/yA+oeLYXXTizXtd7oRb/o5+MGBTnkHHvJUwJKbzQLI6BS9fmZaQ
6Qz75EliV9HbZ0/KSDe87nIw3AdLHJocizM0kZPvNhvHF1gs1VZo8JivBxh/KVPoWXyWizvawkmz
i9Kg8eFsdukUqk2G0Zql+qsOQN4OXtRXcr7r6BtsVZEc2EhRbgNY+vtKJVGivvVIMkTPy+ne1+uQ
pK9zWLcGu02hfPVWea1DTazHr44rTxfnpqnhUXIn7mokYf2bC4hAOo+70Tf0UxOkee/Tms6OoDF+
QVpJ4iUZe9xEvHIGprkGqflaI/NQ5K8HMvJfDjpMNJzppQiYkDoPtmEdz+CkRHuFtnAA25JDS4jB
AMaj3rBX6ANAAAvV9SO2ARE1Upq+MwpgjSoU4793UhvsB4dklQx3FVvlSkbfTP/alV4itQVyQGP1
zck41/fQb8VNW2Rkzd6U+4fo8oIaYc2BX4i7Zd5u9zYmNLziAC84xzbw4DR+fLWTGjb2YBiFKB09
KDbka9D/cB9l0bNSpY5Ptbx79YLwFxJ8cV2RNey15VIeWJdjNS7gyEgqnpEBaiyCyuCTmGp73F3c
5Qlwo7XzvoWLJHk9ePhiKDRd6tODGEG7wury8Fg73R2F0lNNcWkoy0en88YJRQkkcqLrtHTfWLDZ
lGh8minb9hAN0G+EqweK+0VdvPa48DXKw943BLcorvZl7VBPRMtrA8fzaWf3neSrwlAEA1gcmZCr
kY5uK8iQgxXFKpvei4hmmKjJqO5Tmq1EQdXs/VhsrVZycxfkgYc80MsfG30ZX5TEu528jzUsJPQm
wAo4KV3lIiEYMx8xYDSnY3Db1sXtUEx7ni16OHmeBCPgeqMxukpE5rH7CM32BzVxu2mEkroVrGFa
tooR87qFIUtlzJvrKKDD6aJ+44XUlGoj/ysVVRWvywoONajc3IVLtq1TSRo2JLO2ZAWtq31w1F+S
qlQs7SfjZN0jZSDVE6Q5xtT+mRFm9R6l+us/JP3HCIAhTY93zfiJcjgGiKGrOlJv7O+arEyejKKB
HgqhMvCIRQ6FKGRI5izO0zJn6dyNo6+DgfHnpzbYhIFoYjZnyH0kmQ9omudOWkJYoO6ene+mXcDu
ZCiLrsSouUUblmrJNmJhnYTZZhpEsNkD7TYY2xuTtnoJrsDhW1ihkVF9YwqhngGftVnDbOPmPIb+
n0YIYyI/S8/AY+1ei6vvfjH4OLssEbyUfaEwPM7S3kBEQydO5O3rmspjg1bt4Rik3KL28vB6e1ai
uHzJ1ZGqT+78h870QWiRARyyugVvETQ0xs2+8QHt4ZpcnWehWAfNx8VR8oH3BkgEdERlJ2+y68Pe
425pxLtYHtiVEgkFeEw1iyJggRtcrGl1xGQyQhXQtxXqVV7unQcJbkzvW2atMl0ehAxeYdJC+Ccd
2su7djhAxbD98LyNxIWupIEYIFgdJsCjS2wZ4SMHK0rHqnNY069k3JRUmGrD6/U4Dp+6eX33H/xT
TnZsiAqWZjNS7gaIT2yh/Pcrn/7DKSPuNUfIdpDSpbu61sTBGa4XWW+3SyEaQb75BgM4YV2rKOGW
RbivzpckvRT49X9cR2HJThKNsqWduQzPDjEKLagIT45FSQ5D7cGIb3xTn8od2nHnynp92+iSVZlt
249RRKHiQIByepo3jumwQFB26cD6AyJ1YmknG7cZzrs6u2Tgn+nP+VFPN7JBVYfsnjFuzEnqf6OB
wE2ysxD265KAVH8jTOeq0gO8BwqiaT16CQ1ogvjInSl+IGHNV95jmlduHxuVlhqa57bDBhWiw0bM
jSY+PFlxcr6zuXO8ULd/siUiELTGFHhfCaJH4EoLo3NBI9I+T7UAPY6o6vvTZ1ZVJV8EqDRxfoZp
PvO4Ky/bd2oP5ACeH7SF2CUfZrXlY+J12H3kKgV1EaI25tw43p3JtVVj+r5pynnVqyZcskn1iuKN
w4LCUHKxGs/yfRjcJuVaxE+oMuCrGgpZLcemnBXZIHV3leomJN2/P6D9uxKA9bliYER4gaYMnAul
lrNUJ77yREEjUsuq5iZRhCzC14zjT2d4ngSOLHgY5J7ngqES7OJWuLdPtlHog9+yduoGdLlOXBjq
0RsvutzE/5XProCDrLwF0etHylMpXxME3sc5lhhA+7UWP8WfjAvjE8GrcsLIWLIwkwhgrPCeDNs5
lgoadsSDibrEiAIgBgxM/NKk2AABlUsyf4LaB20bjmeMd7jaBj3tcH2OB40HpIo9wrdnqlXZsDqE
G5aIHZKuxqedK/7oKDFgoRRtnKGIgAbf7voD5vmJvzKLmRmZwtjR1Gapiu6nwPjEspxPqRH2mXuH
ZmpAKOfW4FMresBwCN9jM1TVUlEmuyv4lbSv+A9EJeuxZbUyOKJBoN1s/1rZT+ezQAaAhH9ak8hF
auJMsCqCI3jqDUl4bx1gtXv5M8x3ZxyufVyoNOOD9fTXifTG235DSIfjwzgrzxM2EjuIq9rcgz3o
Mb5pYz1neVqxeDVgsbxB2z2qL/ABdY2HDu3f2kOX2WHM8T2G37KhiR117SSn2hIN3vqJ5QevGW5p
Xc0HKvrlc9aAcjoiDwVeGzCzNNbuBCMfb62lqsDxhrm7Cmuql2f2Gu1tKQt0eV9LSrGbTTdkPoDZ
WaebX5Cxiqy+gwrlEy1zezy0uiV5/G0nMZyA8sSM1lrJHob4XiMVF4NmthhZF1CxewunZKmM4i0U
yfSxikQZw5iEcjswv0Tg2DBFZRebxPbyAJ5IT9ehXEAfcn1mJjN3i6UXxvt6FVk7ZSDDmaoCz4r+
QCuMLu61QW7hQGpvQsDqBSeA5qeVyXhFIp89T3KS+/nbfv9EiwXZnzhlTjK9pELKhX5pQ98VvMdp
pzdHc2VtfyfQBACrub+DMxQX8rWZpuRw8SZK4MuQRbyqW+7F3NFJB8r55pmBPBohWypoQJzTrpe9
kXYQkDZvgdYrI0X7u2jxkvNo38aRxWqizFkk2mZW/vKAtV6KH+H1S69nm2Y2ttBIgb2ZfuBf1Zu6
ygYpaSHo9kspsGZVoA92A49+A84t4/OhYtwO/62ujU2j90ykRBcE7rmgWMJhVAPsiokvLYI/cqL9
uFm+5Nnv0D4w0DZuJQdDipHeSieNH/bWqGKWseTPx5uMUYl3oy/C7tOm4KZqgZq54yidYzUEEoC5
YKaFL9EMNtCdc06IKInSbiljXXv9chZEBavctb4ItHkWMbkztPC8HZOmK6tuMbm3RZVBf+2NDvTd
2JY7cWBvtDSgnz5sQStVw1DKYQBS+QHDj/Fyz4cj2WlF2d4pnyHhBG4haxB8IGJcBBHetvKbkdKo
EluyEW55jh8vhzx0TGX8S5IyScVkfExGPuAeZgKbEYd6cUxEUdqj875pFtZkrryC2FWPBWN3Map6
nkBmBXGSi20Hra4flDunIiB8Gv51mDYN8dApbyfvDxhBQ287EmKgfCehjiPJpXSuolY8GVTr80Od
AABWzU41/UvqzOfEImRXzYv2rcbrD4oHBj2QQotA7wL6Nu9rt7C86tjIGoUze4hR4TWgcchVonxS
UfjmE8EMRflHEEEBZWieIoxqxVRcvEj1BWOPpWzSVMQtyRfdmQ0YxiiiNRxpqglUl0MRukfKE7Wi
yxXaI5oEMI1ofpN744EIDmnjD88x+TWeuRYjMSgELM+rmVPKSHCkHsH9kqyZLEKZwl+/qF/avfqr
qs7UbQVguRtvgvpU541Z+SxRi5/EGe4Msu0TkZzG2AdSZ3MxEqxxhGO/WZU8CXyCatO+uhuZ5lfI
3OtShWQoMJAZhCTLiERLOVS+VPF6V4HLI5o0pIjeciNHZeXP/RXoiXaYICCLb/+V4f+9hzUAouzf
Y4zl0MKuk5RtpzfS+9gFpTi06vPqM3Y4kRXN++5+cuhRZg5rSr769/57P4WN4xZYxk6NIWSHB+4I
U6u3AvsBksebaztkprJDuhLnwT+1xm1zSZu6YX9Q+GLLXvnOjmIEadZLelHxZcI+s3gJeb5RGHNr
QWY28x78XoVIBqG9YfbMtl+r2nifviJqV/LVFj/BARrHLroNT6XmD1Lkb3SO57vPo5aUqrvJdM64
A6R72oMafx0VntvUGcpfCUVaBY1BUaXj5tP0o2NUZph1bIJwe1JiWAzpeCQGaKkUSCWN9w2sAGBV
IVt+/vaBEBbGjsXTwy54aB/kG+uG+0objjrHrXX5gKJU5m7+nn0sTk0JUt/pR8q3siM79MNfFNvA
hZvbZEH3xGKsltkmEJyw9yfSNwSLFqX1epQbZYXrjJLuJ5LGB7Z82C6sXQkiGG5M0/iLs72YZAKE
NLeFl/+FTlVWf+NXXMIp88dEcNTvDV2l13zJDeJfgVBnmzoit3TiKRyEQJoshyquC9SZN4i69252
UTWxbXTememfCzGmcy1ljUo9P5CN4aErnVD36A0gyJjak7LCbyp9d3VYdCGMQNErwgjUTq5Cso+x
ur/lHS+YjtDO8+5Gmc/AbwQalf5ntM9Va4aJpMfHHvk9j3/93PBGWe+yUDUKYO4MyRWGjLQPReVz
hC4ZLj0Q2OOYHfAggzUOolpevtPe+mh1lkDeSwJkFkMtDEVlLcP56KnLXLuDD4Yv/pMZeCYTsrif
CJvhnoC4FyjTfSaI0mxFIpvclXw1LkShB0AEmmUEcOJGgS0iTE+1q5Mu9As0O7e9fMGlRczfEOef
VbUovZpQKJWG5JSw/+YDYAtPD8Hp+c8gGyOkcCFdn0ybVaYID3mahN68S1zDk+TJDxU3frI37Br0
BRnlcIL+BQUQh4PvatazxstDqmEcgBc4bt0twZPv503+13DxAiizGoZ+mhnFZUXjyZ1a6J/nxHXA
dFpJhB+mDbt1QRvfrJdxaOxyHmCpSnDuB+j5r9aa2rkRg8W2FuR6WPW2Bs3Eg0f1BxENSPqnvLvQ
xq1oUCBY2oErMR/T4vYPHaYvSGCq/lJdDOTMlzVSZsbxEBOR5YIpz5XJonishzg5hdo6pqxxl2yl
ljOGe3copPi9X9rD53lgmUI9if8lL1H5oW1hFFtznCbroVPyTT57xnqEhfwtLEqeNse+RDUwBAep
IFsBGKvVTTZua/0svWuUtgU8b0vPRBfL60xqRw50GJ+nwzq5nC5o0IcaapHvuiEqjNUsvF0gTqz/
L2fOulrH3A97g7wGV2YK/W0EFBDpO85iAz5keksnxfGot6ZJ3AR9D0iJUQTJl/uEj7q3k2cwWUsM
1DtJ/0iENd6IQtUiE7oFB0Yitj2Md7BaAG3i1OW216Qo6XdgO47/u9k94h/X35ALlbXayWeabXZM
e2Rm8yqpXvF5+hk9IjpY3tQfraMGL3TGx4EJWZh/yuEXfMnQHqhnvWhFuoJT03dmAQO24PJ9sTQK
/LPc6+Q4JaymoPX+Sfc16tgifJqsx2LPwwmjBLW4KkYilgCvlzS+a2F8x0Rue5Izn7Lli8ad8Dsj
GDk0sS66Qym5AGYBbGRnS/PP/zjsRRx8M94lcQ5/gY7TGddOhkQlwvAEG7KPohlBauTcPvGtg2xc
Y5K89rvUSrlB44Sav31gWsqn5w3AvegScsAXnYZzqCKMhltY3LocjNRZO63vKBZX8tCIBu1VDi6o
SQgH1DON56XBdjzgDa24o7q8fKVF30OfKcVy8TXqugjgF2IpOcnL/P2HiEcNzQ1L0PZztVQ2NoRr
VSQfeWu6h+PxcEIRj8aryfW78FDE1uX1OgCDkO/VrruNNOvUSmD0ICPyqDVWw1KLg37EV5I/6ne5
23sG9uC22kOXrRKAG2wowvNvXJrDhX+fRV6fexzZ3Qfge6VLp1mU7jlm6xNXb7hD9frfyy8zRZrS
C64WFgKuFwbUpIhrLiskGpsX5AMACjKMd8MFZQ2iRQ1Yfn8G79Sf9L1f/T2lZSAGa1+8mY2uAMpK
wLDqPQZIxJRFMqf5OrZZyl46qwjBuhqShGTdRRmc95+Z+MXP63muWhcoboeHSEHWhdv751Pu8Ya/
M3yy0OfzzJnXPbEqY6ryjTG365SMWog2K/UjadXY8arVYlyFeE/51+DFQ7WRZXF7FevVPKoCEM5j
9wxa0cQIAXJnHfrqwfEj4KWQrrDrSqV/5AvGBE/CzVJAngi9r/3HRYHEYIEppcI7Wwh+reXdNrJG
ygzHSo2q2YyHdwhrNfXPEpcWJYdH/Ty5cQotKmDH0OIg1KD9FtKf0I+t8XtJuAPUN/zvQuJ4USmD
zWRr/bq3pL2x90vk9nMnJfp9SA+wSlEe9e1zlPB5+ad3uBBvbgyPO13y2RHS95nh8y578nqEuaQf
GdsuxNoNeJnlsnH2azfZeBJrC37Q/1b1OTBj/xlok8rZ2yqrmDP8wD96RKX6HyH2kszjprd6DG3R
j0U1jqWvgtJ+vNVAqt4XmbGzGToJjHpVXYizIjv4YUO+QhDrSrAYebp5ONxA2sPMqtB41FEduxkG
psktgj4ZUAd6yLjPBPC9LOTwOMTAjPTtboj6cUnH5NcCAi1uA6FsfzuQt6sEFiBkonYQzfGJGKqT
ppW0W+wOYNVbsT9/NT6tlqhLb40rGC/SQvY9I6F86yr9um/mZWIQlPs5q2eMGrkdxUG/YOg3VvUd
TRIkmaW85bORkAMsqT0MR6lzGau5HU7ehqt83s+DYUFIB0dZiU3Q3/eoIfG9w/TBeH7HQJZAGhlH
NeEsSUwYrTzAaQGVwsZaJzpiJXoWHHY2J0TcXXXqxAqxpf1MS7iEAaSso8p9HMyhWGEnO904gnZy
SUzjWzkvJO1CCIG5tPAnIss1FwHqzTHY9B38byxMoNeckSKNoXdZJYYNMHkC7GBBxRczfHpUFlO0
rl4elVA7LRjR9c7VLV8P5TPDv11Wzww5jxbT5bTXEj/MGu811ziK3cnUkh5fAEbXVMrV2m/2Az3t
34vHt1RFvPpg0yd5FvU/m3qPSXlFLT9gVY/ntxLglHrXKrBO2+4u2+HbNYUYFgnTBLTyy6fCPggH
+woztysuG/pfeEbxhpEXOHeUot6Y3t5ttXU/MSP0Z2RDMJiHm+h54v00omjKdG0vuXscpxHp0ahY
++5dSg4jzxrvCqMJO0mANfuLp+WLyLptg0hMO2620UalZKh79kmf3qiuh86FqWMs2yldm93XKqD2
OeQiwiT4A1zIyl0q+15RVvfX7F584sQ/uLLEVcJS3aMLt1Gd3ZOY6gPEVe4YEpWG8aaUtA7AovUR
3XYiB3TW+aFoMMneNoNNud/3GfxcbNKxH/+V7Neo1IeicF8EqI9MBRsmehZaVOq0Adrx4e8hlYX+
Zx/V+54jPWBu/cnvKtoLjAzg3yw7Su+KYVGFsEdPQp08qVF1dE0rjHhkDCCbKPKgi3zbeT09hi64
PFfvQfD9IqWmB9hVBUHDbtyUP/L7s8CiO1hjyFrFqty5ErMGFjgq0l9cUC/V0Zk0YIjpwyOP2Enc
tZ+bZk5Wp5eyJ8+dA5SaTEg9P/6ivIBD1DnNPFJWP7mNjBbdCDah81V9GTv0cFZkHN37NREvrkbt
2ZKqD3bUBnywJZsR/pp9yL9eErCFQiuQm7Ximnd7ofqRr9+dhKhe9B4G7t31eAQt5sOUJjikIvHO
JAaX0jk6kJ0W2ducTT+eOryWd+OwAzq3XeDwOItx0wd+qSmHuDPOxRHb5IOGqoTzGADMkGsLNKto
x/kYrySEizYKNGl4/mQkx+fhZ50N/mRYmJabMZAOb9myBpiHEgTpS0ZLH0NqPqIB5C9UfKhbShU+
uzOOD3llYdOtRIT7iaVVVHz/drhKqENFMy6C7CFZdHU2Kt1h9Xwz8o9HJlrFs4xHBi0wX2l8/NGt
0hf8zoDGEOfQUJGYWmALG3jTsKd6HBqCoAJZWDRGF9TDCXA6Zsam1v4H9wl2spWuD540i0aPvgf1
ZEgf8775gEdXGTfbR74UlMc6B/UqoSVq0LmO+bMPJlUPUvL+2nGN8tKoFEeCyMd+L5rZ2Z0+pf0q
XX2/E/PXk/XGzYZZK4U23NWUj8b7R2CgrSCIV9r8/J5vGcWGjfS/8wFVAmSarIC0qdjnKwpX69e6
RXVHbTPyK45kR2A+H24dGUHlRcVa0IK+zXfg0IzaK4vaN/vfPyno/ba98SV5OGo/7FPrk2X2HnMe
3yPYBjo8J0q10e0UN4lCD0dB20Q9FW67lnMiPWVuabwUYtnox07gtf1Cy7QVFdfMKRHjEsRSxqtC
aNeH7INHGF6IBXDN4ufNUtRMFrt5dkEYY8DKUTfuZe5YWLCw4PnIQkhk5A4+hIHYgKunQxdVooW5
n2hG32r89eJSNBcCn33xbkKSmT5nFwgfiVw++BCM+CCOkxNODnrWfVgNUtf38FAHs0AXs/J9cwcd
s5nHVfjnzpKDj+uEm8USgFPY8VXiCCj3/qRqnjaVaDIYD4bs5SXCNAOo5evTPPxmXrdPvAk9jNU6
LdD1NV/zT1TtCw5LrTSPQdLBcvuY3UaeIf+BcJQvKDLc5h+z5tYsm6I/cUMG0rwIpQ6AUa8QaQlJ
4bUilVJbw12BkgoGOOlrtnPIyV0xME/t9XT7ohqhBZg0xe+eyeUp/O8AY0yM9Zp+c5G2gLDNNMlc
ckdMwVyEy8FDreD0ayICgEpFNcAelglM2ZVwRjm5SJhE1r+NQGyl0lWWGqw3532ocemqwwogVMvv
O6sm0Wyw8ROFIb2vaDrkufqjiVPhPcWeBklArboZapuijnqJC/i2oo+/kNH6efPmDY5Lqbm60QZp
lBkBmiBmRySzO7JPGcXJ9WuMCR6ZF61CbBdf6t+ZWFibGo9iokP4CSxE3r3NpGI6UtyGEV+RgQb1
YPdxafaqZYjaytrNXPnB459PrvuR2YTaPQL6IvoYLusK+tHxCDDPeTKBulN+q+bLO2egxAaGSXUh
8+lTExhPKmeeBhlWYzABLD7HGLk5cpleuMl7Vlmfr0icgsht48kaHKa2rvWfCrTU3FGBl2Z43piy
t2EN9/wvfsrB4GT/3hYczWHwMXFEbrEx8rbKtupziHBIgamp7pS4uieSqL0rGSNsaNk8L20yw9zS
Vt9tjlvg2LRFcmtN/LGVn5Z5sn67K/TPjbPaFMUNvfppqxTyXHrmn843skOC9Rn9LaF2KglpocAX
lnJua261Pd/yYQjL+kQ6GvI9M6IENsg6Dl6F7Pb+Y1cvW0LT6O93Z4Y30+MFMLS1SbvoR3/Ci9nE
6wGBZCJe4BDg8sXKwcYK526r4Tiwct+j4Qud4LVeOixBCsnspqPKLoYtHFxvPmRAKSi4/PBN9Klc
VzV/Xvvyo4KWAV6rZYc1qqQyjqhFXzSkkDuIJ7Okmp0Hty6TkbOEZFQq+KLGPD3yURQ3v+rrUXkQ
peIJN/JKPcD7xMwbnRUMBBtoxGpo9TJf5CjB24GW/pAr5NhUYNejl9Vzj0ItSj3/RW+d2eG9Xzcc
+H7vu/FF+9GT+Ek0c5Ej6IEBGn/AxF4BqmL/+HR8Epn3FzmhjnEqzzEJ7dv70SEIzW9rGe2sw4yD
0Irxs3eBEc9oAbSiLqYem7wl9puaWpyrzUPH9xNXRvjNDLrgHbVqwZw56Oa3pH/XlS0OHtKRR//y
zPGDQGAB3uOLAWDkmvu2uXFODYt4lZ9yhklUuzYV4vIpEgmMR0qcLbZXUvOxoeF240VrNzPYBNVn
Qt1wqfVQCuQxoKxbf5c5XGdDA8KwX+wCiaSOjRv8Jfuw5E27HI541gJuQjcTtYTelSHs1Mvz3YmU
iQGw5LxcBYBnQbCI2a2QByeaVV85MEMPHi7EOo9Nn5jzHPkJEULJLWBRyQ1/9KTIYZ6WcNNrU7Zg
8+z8ye1Pwcb2TYaN3mLhpwNvM9hrciK6QPlum0InA0UbDKbF5KKsxHaQp4Cs0qrZXzo61h0dfoPt
C0DKzu/k0ojCmnUtffpwuj8vhwIUtjwef8+/qMpXHY9ghCh74PMBQXwFTtwdMcMjBaHOGuO+S3PE
n6eAOKeyMVo3UGHz4Fb6G1vG3YcRvPF28Qm5P3yvWJh+IjOWdWxMZcs00AAKottiMxhnNacLENaO
BJJKF2PI9d5LpGhJfZ6l6KVFFeP/SAZu3P6sAmqPh56Gk6lV73ner6LGVRRBls0XvfiWamaKYXMD
jl8C/BDRLjLcNnKKy1Ye2dVz/dFzi45E2QPb/AwDlny6gRPBr6rVIjsv6ic87nw4+Vjj/j2zB57r
Lnbt/jykZRsC/boaBMCAO7iP5pP1LN9BIqFu4VkVdZhqKg25GjnYGAMLmlEr47r9FWJLv91cXfh4
1lx+VCUkqvK1mh4gvzmeWRVmVyQv/hxgfZZdg0heCdluidAH4Ffdn9tGGKHiT+untk7FXjykOei6
Y5SSZd+UpA3JwN8DdwuxC474Ys2WJICl/AArg+h5ytoggI534LSKNKDV7+DHNhPP6pciw7hQg58I
sY/CpT42HJFI8Alu1JeQVOKnTIoksJ4V4r4zcIWp8U0H7hnpgREJwpoXEZY2NtZgGKx2cS9OR7aB
Pm2Zz8LA6hqEXejiyt0lVlXqwYrxyUwRFimsbS1pn9XqZATusppUNfjW3edODzodiW9s6XawmtOA
NbGD1HZv6Ax7PPTXkkXXdP0QxiAn0Gz3qYJ8hurMvYZqeMDe8L8vUldDxuBnuoTQCNlMYZZ9kAj0
z2rKQ8+SLNAfZmd+VveNRBGk2EZ47FEopSQLeYF8eRxysY1lSLubQgnz/MBsxxfdES+El7xll5wq
HcnwIj9uaUwgjn4oWbWGlJ9xCeZlIBFp/e6zLlqr5IAQCNwXZHoOAVavybQOQXoiM12dQDMHmw8t
VTN80IekUiP/MYs7yQxol+DjRyG3+JbaD+X4p0xxODGYar3ltJKBlFLuWHfpD/a55l7T48yyPYwa
NpSLJC9+0ix0OSpFiuLgIEBGE0LKUjbuHtH6YI7ygipGbGUVjPuqrSzJFJ08uZKkMR8HT4bU6GTj
Xe6X0S5iLhoAiEZGNWXNpgqw2nCWp9dKgH6jgOqsNk92qjL7AtYZyrxB8rCPEgTJk6bc8wQzH6Fx
t+wbLUs8+CfL0ESJjKnei0A2Np/pirxVy7xVkyiqR4sR+a4H1N1SwvpoN7NbjB4IQPjxY+TKheEg
3iyTbHy4GDdTWrhjRwr9JHEYrhFjpvyLk8+H8DR1JvFwMubD+IjeweDg9VZ/pSnI01a9+TBWXBqa
ak9l0S8ud4Edbex5RQPOHJ82FtHMWssAEJP2VYifBz/X6jn2cs0wneBK8ZUIJUPNSNIDjDWnCxUM
UqC99itxej3G4QO+51L3ghAgxIijkEqn7/NtqpmElvomcO5NU3nEIWXHT725ndsU9y+5CXwMKguW
MW3RdGtWzD3RKq5xWxQu1eUJR/p/QmqzTE+g2BBQcF7ouse93OPNAvSnVkoUb2ufui7eGcm/23w6
hleUerjp+NdifnrwjkAPBfWx9c0oJe7/ytj2SSJtS7Xz/ezca+RoFbo0W7xbJfeCtiO/IqarAAoj
Zz0F869VrNJdtdJlbptxzr+bK2zTNM5zvzPIcAR2WFWP3WcmvC9fUbd1YUl5BietWAIRC6v8gGY9
iSUhnR85ccoeNPb+HxDcqbZm2G6u/FXfcATAKsNHVPFZsIqfewdSkWskXpOBnmBFRdqesLGdjuD+
U4+moZgz17E7ZC2EKC8du9dUE6TZeiWpv3hPBJiC0mXQ1Tssb0T0ukRoHWSqrBlex7BitxOgIqK2
b0SK0nNRTUV7SptrdxwWND97gWYZ7oOt3neS4dFO4R/KY6U0Cm3CtFhU2kzDf61qsKOB7QiI94V5
/VtM++gfi6TLdw1dLgDd65eZfcQ7E8vpY7QzrmuX+AWttX9ZaT/ESBxhViyDCLx1jZ2IaNwo8gSG
CCPAxRQZPZfPNuM7zm0Cz/aFJA1kFsgTH51WS96OVqAKusUccJkh0y+Q8s+gSC6suLhH66L3lPeR
bZf1Yi1WCeWPUv9Og8oHmVcrCqyqAGeJrK3o3IIRP7A412ExvAyAYCS3eof5eOp9qOVmzoisWWV5
9D+DUsXR4aVoHcqXjECS29oWV/g/0ei0lHtfFuUywwtfdCCWAVkipTS8ChAy4qz8Ek8uSaTArlB8
rktKnX/LW7q5fKBhwkCznG9BHBHJ8K4tlEiACU4UrgFw2y7UE/Ni69pa5plXjbPTSKPhHQJQp8yH
lN7jXE7E81XfUw3fn79IVPks4vzt1rRps1nL47s7zUH1LQfEteAe+snY66ivrcRb/61OJUErSb+g
5LaDKXhl5p2G9nacqvW/ohv/oipiu2ClPyGh+pnMDvo/PCdR+LANbkxeEkjUy7rM99czlr9oMxZA
kC5/D6f8j0rbL8cXulweu/Lt2GKNHQ24VddPyZPkSpwYUDPktO0UFyoCEDqueF1749dLEgmH08cr
0uzu1bri+gpzFcvzH6kfi8N0AZVs4TbDPKIU1pstSrYFxl0sxiJopfSAwX8h3dXwJpiZrziIvT47
xbanMOtEscKRMNStc1R3Ka6iXnexEk27/7yOvrahFDjLC+Vo+BbMdTbRk2LX1c0GOgq0IzfYdLDu
IYEwMAlQs4CLFO6/nsoPCkQr8e4JhiMy1t0IdElUVjyho69se/zRO4GoVrMlMEOunwdI+VKBtIGd
760a4cUPL4Hn2CLtSlIsWbPCRBKHoY/i9rITBrTQ9ez74sisNTW5SFOd2bV/Ji9mVDDK/qeX43bC
TzmFgqTQEsi5P0vb9cokVF5LBQ9qjCvw2u2amrwlW1XaES60BK9PplZQ6/MYu8dTz6QqS2eH1MKT
+BrmP8n6AJkTYd4ijMVhau+LiKeEGyD1+sWGrhLtYSaFXEHH91JlA4zyzppaoUqBnY/bj9Ir34kc
5OM6iaKIwkZBCIsG/i2+Dul0bCMVmAAxAW74QmkDUwS4I9BK3UpnGDFLKtNjmSxmfyOKF40/51fZ
JjnC/6eSX9PPJvD57TzhTX9wWdhiY18+VtwoNc9YLCyfvGeyXEyLicwG9Hu/wI/2whMHiQXKPBc2
1nZNAYYfYzLjVcf7PaI0ux6de0Oh3kX+7gvJ6WXe/KiC6ekVN/aYvdN4cUEc+YQuftfVZ1/LwCSE
Jz5FPIiW7ANgNabFXxMBFvUG10LyIVdDZJYHJQCYDO7yfO26FFU+9vww2si3s4Js11e5QiI28F0r
TGEZa8YynS7kZn7UQaUEGl19PUu2JnUZeNNYq963X+BIVgfbFflgKnHsozRV89mWrWxmkv6dBR02
K2VDcuhuDQM/NNObT+xrkZASqmTq/Gc/yCITir+TvPBLB0tW7D28Ji5vra4zHHY9AR5r3RplHBMh
/wxZG4aqT62cmL4gBgbr/aRAQfdTtLerYjcEgTl9h1DR2SSrnN47Vpr0FNb6RGw0a+Yuyku2mR0N
Uq2CFVKTh10Kga/xmjjEtNV1agRSfefrTgeffkBb+kiAk1QU8poSKLZG57Jr4acJI0ApCmpAS5eZ
2gFR+r/shpfBFno7G3tqV6lwgWpkgFprN9+lRD33mHkdkptFscDv48j5mhjmlHW0g3MsMTUjkRDO
ME54p4HVQzgrT7Cd5ShFQ4orpbbKb671GhUtQljAwxU/kRl2dG6f+FC+XqAJpPIrUL7p/FnYiBnF
nRfUp5JBtUuWBbT06y0ZflFZmUMihYhuY1SRA8pKLPpXyRO6O8Tn2InvZRIk2Yy3J4zv17senAtK
KSn2bfmOxmm64Za2+K8SWqPKT6DeJCwtyNF4huqU5e6GX1I9E9tVNS0bRSHorqZ/NSM32OzbuGvV
9BCTR9OxW6fWXBFmU5vzptQbTGF1D7NyuVoyBsLmPOY3VNbuf+iOplzOzT/RqzfUvuyLZ9jZXhj2
ACg3g9YHFr4vrnEGQgk1W5qfyoa0LZ/5it5pdtL3jTSlx2WHbUDl3dDfh2S8x7e0CeJq782Z2Lea
Tz8d+rl7vl9sti/dNpZsKsnGjoRb2ptmIH32cF8bVDO6TPp2nEzS3v70X2n/9D27lg2wq+Q6b1q8
+kzeUdmwe7zlBwb047Y0lKczKq4yv2ERA1UfWEM2CaD+ZBlYeJqcp3j02pzBj1yBNkTlwp7QglEF
k/wc2qattDJE2ThSDOGyfxnktt8/3S1YRF2nDiE5fTXPMFiy9NaJeDBnZBz0/GXSOQsNaYV8gAms
oBbnuWcnXE9VW/KifGj4vs1qbGbQ9cRi2ic4F7oTf+TUtFgHs3damIwk0xzeTz0Tj5FymWJkkIpw
mUdluwJN+4JQNZ5JJfGG2VLbJIuBQQmHw+8RhkvrEx5xd5huA9bFQHFK9J+D4g/oQjOXND+aKLMb
UPLYZECcZBZyUhN65gUNIEBDT0+uh6/XOLUqjY2uy9QogwscwxcKE0DCk7PTxTQvut2knwd6Aj33
Md5pNzRg5ZNHrW9HsGPbolW5QZ8mZK6Jm1RcGABZimy01RVatKDR1WXrDqMr73pWMlU6MIaEDj1g
k3+EvIwceNWPvqaW5XJoY2K1yRJHQzuf2Sz1uHlfUFNIhDWam81OpfzkIZTDrQRamlcnwKeP0H2y
7wDiTIi6Ixru2cbcOgilt4vXuZt1V8Ow/6x55YB0m8QznGr3HUyD9AKhryGXy7tJbUUBQMiIT8yb
Lx1FMO/9n7wBX+9LfIRuP3jdT+iMmr6pbpHaESmoTqrgkC0HkfyjbqDGypW49zmK0lGpLYEWkjB4
GaaDvuQFsJ5nxS7v75Eb+lwYkKsQTTOvY5hJ+EzDaZiQ8D3kQhEWybZgE1KeW2ah9r/k8SkSA4eN
R3QV5t58h4UJKsJGjSEjPFPAN3BDx6V5VRxb6s8pKf0JMUykdteYgVWsYr66Y/Xr87ngkTDROQ30
qYCDVdN0A4TXoGfhIwURnm8ZeApzluHW+GmdG3srL9vNSSZ8MVrjWvE28fmU2Zk6DTxhxEf8lA81
Qafq3SDFaxVNBtOtuHTBpeqgLn0Vj6sAEaY792FKhqPW9jfESzi3XuTAtl0CvC4z/Z5v2TruxkpQ
iavp1ZwuQOLlap7665dsIfTKXLWfyFbXOC80eTPO04tjuGnU8KIzQkQ5w2BHK//4c3/OdSZwSoQI
7MuLveum2dHnOImofLr5zGlsuSZrh5AauX6wwJGrvsGM0qqaedfxXQEBIzKSuUPj1eHLnMZ/PZZh
fAO/r+u6cgsOTj6OONbc6ewvOk4hTVyYzOpG2hsenNElUHYD2/ok8PCT6bDpPhcmsQoW44xicw5A
4Bpupk2tB3oA1XcfOHcJ2IgzHUntxqRq71JHrCOtB0wq2S3TibekSjsjYXHYMVw5od250YgcsZXW
CmG6VzNu1lk4z8QCalfvRSQM29H2XQa9CaXjG+EEcf/0F+qK0/sxmf/e6EaSP2ljS4mHBepeWiKa
NFcYeQHPS8SGRRi92JH7VJdjyEjUWSPGxM4qw6IC0bj4QSXWU+E7MjOVaTxixDduHhgKasZv4HUO
2LFwZxtZM+BaQBHIhW3agT62k1ah441Tn5HkiEJgUKxwGFi3bDtVmq+izfWdu7JL4rxkF6TXbPlC
RehWy1gAFzk3RogEIc2tE8cyRJNO41OwlmsKz/yvZbykC0bbdwjIvadoNLFUpppoH6zHf5evsprB
1fzhYA9ic+bQWGgozploPXOYnWTI0kIEZNf407sdpAKcb36j8tjL2Y07pR/N+C7AGy7symNAg6D1
Tmn0OQTNjqZtMfbnPpWhxBXA57pVWa5SnOlxCzPyHV2haN5TZHRNDAjbEN49giRLJTcaLAwsI+57
AGeQ9CVO/rmMlTwsFEq2MrrGZVygcHl9nhbAr5GRYtbo07eL+dB2tCXkW3SrbLbofu6A9VUL5oLd
dKDXsFIwzLlt87/yjBdo26TptWxElvj9kDXazC388wKrtx6JCh8tEgPlGrSAfhHQYSp45s1x3rn7
L0xyfbxwUmBcL6IDq6Scl1Gzf+rCxM0tG4pFR2rXoK1jQYK5GJH/f9XFDMpN15nMiUwN4cNBkaWq
ZYyJtZgbSqDS7Ohd2f1E0HNkpMfla7Wjb6CNjMNZH/nzPs0ZH4A7YnBNLtg/2f0PilEgL+xBYCY6
+ESEisEioeliYYov5P/+Vi5W5R9HkR7aSNwr9AHrxLoo9tpkO9MvP/4pUhiHdzqa4SL31PeVHNug
8PepfOjIBOzycnAdZ8eWZg12vHLAUtK0IP/FJ7bjrT4ghvfCZTLitwGWO2drUDUeekkBT/b1sJM4
Xe0qR0AoJlWNYn3OG68d00daRGFRSKGk/kU7kqJYJRplloh55Cd5AyZLSWnzkjSjJ0v5DkyX2k9z
yz3Oc0Z82TsDMtuT8usz7PulTi+f27xKih2LHtjXD1TOPco4KkcLRzC40R4QCgQ4c7XY89M9bmRy
WqVE1qX6KZfYPevP/3/HtbwtMJQVEYfP7f9RHzvcJZ/jTacD2kXceOo9driINGlpRUJOluTpplxL
AP7ZjjQl9eP0tcImuAK7PMtjIlQtgcDPlaUPJQVHBgGY6eaIqUDtxyLxA1DPdNk5i6TjBal5Aahe
obZboJ5pf1KYScVvGdP28yPdI/BXp/V/sKTG4/1KCnznwf1CEPgI83HAPCvY3Yl+jclALlroCEVQ
vzBDuVfsq0RpbKXfNWkh9K1eIpY87HAEpn0Bu5/6Qc8lHNgywfW2qPZ1B2x6CG89r3ojRD4HpQOQ
ryypvRW3srLRYY9M24/HzHuQrz82AKTFlfAHYZZMcCMPfh1Ue0J8C4tIxGY2qYAPxCiYJf46nnVi
YJRmsm3+PvaXnwIOBCztMDEVAhhKfZ8jIGEnFSXHerFVBgMa84v38L2HjKymq7jzDbmkD9OuRFl/
6zCbE0DHaZR4PHXT9Lv9o+w16uwAp0l4aUKC08SGbWoP05jUqNjAt60h+t5QOVtGsQ04sT34Lc+a
pXwIOrKtHm0+pXieUWV8eQhT6OeZOowucgIkvtLmQnAN+K+PEPzlGLJghkDm4aDIUqgek1pXvQhR
jiPx/g5laMiWXu9+RMAy7zW7TRoWNj9bdv488KEvR2hT7ad+ejoCwh61WgGxV96pvdVo3WfiXF1Q
5imXGt4Se7mgnZoEpxEQ0vaMzZv1pN3nUndGNnfV8I2+0jh75P2UNjQT2O/VyCD+//Iq4zFW6LuI
XT59DP+6YFQ/Uu91PcBT7us7pat1rY8yWwmohiHMAwcxAPl7rK9GVuDbV1g17W/oxg8XFi0tna9e
MglKZgzBEmhxP3xWwtiblA+VSGlGgNcxgrUYauelmy47zRPpXXgnA55JEwIfC70RCmCXT4WXJ9H5
XEe0OYrcmSHimw148X0L5hpfsdU6A6lHw8zHS94UzB8Be/osLx2RocZyCIqL8KgOFy3XL14SxPK2
IBqrOVl6emfVxqtp8C/tY3o9VRXVfAhuonKy5sYf0lPl7KFgMx6CxYijY+7e7MVIelhJtQ93e1YD
oU7CnOwLe/TdywZZWka1On8MwiVl5w74vsckC+s1nRW4P350Mowsi6ZasHwXuiSkGnmEUpiHZGHl
QspDrsuVu3YXEwD2LOkDbqVDalinfX9bFc8B1n+WemdlLVwIORByWiW0QgbqU2QUhhWmyFk504xL
/l2iMkAH6UwW/AEKIsL1eZXEfX6zjs0GsKu1k02qWRYVSsC4biMNmsVAZjzQm3f1xLh8U4VwGptp
Q8Fv+7f9Hb8RfZVjeiAXedLtENCG7TlA6IOB7xU+SYPTD8Ido2Vzc6EQfrEYZTxR64RF9BSsBKB5
Akd8lN0rBnbFYTlWjlHiNISrNghv3wvRFa/cYKfDQpzpm4pvcFX86ZZ41x2w7OAIUezagMbl+J+3
bsj0ez0IsEXHevaGGZnx1o6I8tCJuoO2vai9eoODgWQxN/1XoculZLwPmHGz7DxS08A4YucCYl3Z
HXWv9VEkWGNZ/VlG0JdEBUMfuNedA8/UFrkHdRUzGqubLKMVVFF55rwenvFTrpns3hzeVQAIMXWa
GGm2VmBuPOI/96dEBlND4tCTa5DM7nKhjNOY/wyTCVMmc82lUbrjKvV4iRyORx/Tw7p/gHKKKJ4M
bqfAUwg8qNjxmOwLfHZtL/STInl1J3bxq3l/mdOIsV+mmyMuJ7sr9+woe5gyyE05Y8YmPxozsmaP
w5JXa+ezFFbt/z5Sdy4lzn3xxNlRqNJCNzCFHHaeztq8vgT7F1EceUeFYEHOOCWB3kQjFmGEfCrO
WfYB/Y+0ldV5WwihMDwJbjIKh41mMklk79qF6oAmLVKYTtipn9QwFzi8G451Nd0u0Nu9oDtEH1Oi
+kKPYVEbnGDTRWUG0P2KgaBZQg4vv05kgQMK60u15GbdIZPmVEqnS36FzzfV9SHDX3NTqbd7qbEQ
qnPPVyr11UFv3XMaor+s0XD8luc8XbfjvgqnGf8yJYJeU+rKPxv1mgR9Jv3tsZ8k3BoiIAH1HgXR
+frKhSw5nSFGaZ20F5BJebAPY0arvObbIPz5TxDrxZ8Ib2oNVRKFSroFjRwHmevixxXnQVH/dG8P
0UgH3ulQBs3Tu3Dsd/jJGPWfBq/QzLktszCnbEPQEdybtFvwiCUTp3b/ixn43ZqkiBf1wWK9d/aH
LhhrSqDC0I1oLM/RRmV6kBa7sWJfJjYMGuf7+Q4MPLCdaY3m/q9lgeX/Ph+CazA8dnE3Zk9gcxvv
999FCecvjB78SAWpnXUXOwX5KhRztmz/7fVfaFI/d94NfW2zHDtY1F648H2E54jS5CoYtDoIqde0
eiTflH86d0kEw28Lm5Gcp1fQt46wd/3Y36Dh3T9AksfdtAXKRgGWV0n2nTGl+tGpkc970Js4+jU3
dPs1dglmZHrzsmIOQzC16QAYMAZgxl237sMf6zxYtz0zR5NsGcH6ri3ziDjjWnzNasXY+UIwZdto
ijnIKDuqDCXz4ViG/FmmvDshum1wcRsTaxicq1zFYqAxyDCLsA7FXB5rz84IXgtSVlDZIgWrlgpv
P4TrSt6/hvlmAZ4s1jvArMtA4TpLj0eKZndzyOoLq5m81ghgWdSQrfE8n6TLnsKK1UVnTaqY4fuU
3OSHvLaDEe09iQF70nxQe41LDVT0OfuhXPbknP8d3jSdypbsWQLJWxW6Z+n08+VOisUK3fpT4tdX
DVb5PlYulAvbXYFXwKTYpU1HM1BzztluK96cSqTDxTD+4pQMxoq6aaje7AiFbKFKyf7wJi7ikgSe
z0niGjWljucMKKqHcmdR6XxQhwhEJUPtPHJWWpyMDqUnrBMVtICsLMqpwDvXU1gQ9UhcwfLXXWdo
bmd9U499kVGc/RzAuCkjeQ1/B609umtzruxaXsoy+yZhwAAftkDoSJeGrEdvHPrRz+hydiEtl4rZ
6Ky9fdmLWkZKVryZO3aJzfxdFbTowuIrXuaPglxvM41hVwy2ruDM+87O9Rw250Ew2iWNFt9w59aa
SPwYJi4qqY1WLDD75sXmhhlqGou5xCvfsPGTyHWaX0li8Dd3+EQuHTj+B2LH8vIVrlgSBlPxtVY7
PxnWmJWgeGYG8u8yhNsm12W1tI0M0D+96IrOa6ZbTpRhI0E2PYMgii6+1r8dQtp3wXvAaJZ+Qp/E
7oNCSgvZ76dgVNq6zIINMEPAdZlVX7D2INXm2wlcMsg6RC23AbyJmAuhELi/Tle2dOg1z8xLgVQx
X5d6FhwJtyqQoH/g1YuAPLcM81jBpKsFmEo32A7lP7yRkTYy5K7JwKub5hThTztDXjWsvyUO4ked
9qSH47W0m8zK8Amlp0DEXkEGEYPKTGZGpg/D1E/xVWEBEdsPJt1vyVXid45fwE5iUc5ofC3xp1+1
0vSfDgwKCn8sOKeDIdcayCh5EjddYUWH6wuiYBqkET8htKbEMJ5utH4tCMTcuhYWC6vELyIlTrHA
TBS9KAGndVvJC9mEcr7PKGHbu6PpGgBRVqvrquL97rhizC9pPr1WgglxB2NNLi6SiSPlCjBVDYHJ
0e+oQknZZ/VAn6Y6fuHarYZsL/+DbyWIxefRWSwzkyBMsIAn8fy37rCcWeeylRJGubmcmK4h4lnj
SWl7LsRKFY3sRdWMeeoS4lDdwTSCs1Y2pKza3zoCXnUKL42gKX7GAqiYfx72ewx0WDlXi+d3YR1/
R7d94h3ZYOmGCfBC8Fz03ETtBp3PTCpAAz68llDcuVHCH7g848ehYYlDuI5deKXGSnMGdHFJdAj+
9HZmSMBT7hcNQOYjt1nfcs8VbbHANvd43YMei8Rm9vQ+hcH/qY6ybevH9ZExCcdbfezJ6kGD66Dp
Tu+Ga6yFxvlxw1P62YM/wJIiOLmaB8+hryroujRpgpT+7sfVUdMTGmDTOYvXUMEXLW2XaD5dRtmB
2LwWUlLzeAvVTTSAeDN+SnVJA381sNpmSuWvX+nwQ2YnhBovTM7v/ZPksAt8uulrD0Qd54uwuOFM
Ts/EigFt+nLe6SsQSArk8BgBlw/c2z7239aGeF3E60EdP8TcLbGYHjSWv+LKypHh3P039xaTDLSI
NuI9Tgni5KDus7BRuOP7X1NwDD/gz2T+xdOlUVb+QyXc6Arjg523H+kdoA016rHfKf6wz43tLbMo
LQDVGk3n1X0CHKSOXs2cA0I2vDY0CBlYiJV5yxpTLndfKV/XKRZCz8LuImqcGUn9HbIcYoLLOwSn
iYaQRANjlzTv5mPdGnp2pHBxrgDe6f1/EajMD8RDBhRYmVfRhePQqGVkYN3KuqG5vb9FpGcZMgQb
gQUNQ68Rf6Y5u8MFYUhYuP04z//Cm+a5tLnhIGegVTakYJm+04mpfTkYj7opfKfC75nR4Ai3xlMT
SCQBemglzZxpJA7zI4Bosl/LgmKGziHM8g4o2Ctc4J45dA0vDApTKRvSCmtAcVpBPpdfdK0kqs1B
2yHTJ+P48HCJQvFhFqtXlkJYEjnLkhCCebg5gr+qd57FD85YWYH3vGOJDyUwAKqsVnop6R9+JteZ
iN/GpDtqmMMh6+M1AEiF/MuScBu6cB2LNch+tVS14Us2mAT+lgDbsrGJerqu1LTYABfwatGWQLNj
joyCb6ZjyEBSoitOnvvgOq5InIj1tb6XitvHnbxo6mJ6U4kuR3D4sLU3xaLvr3oMKJ1Bi+XUhNI4
KmmZHei3rf4mC0tapO/TjEMY6KQ4+KOTF/xoPJ3QtZa3skYXJfpHQX08/KwoOoo/CJt/vONoqh33
PYHfYGNeXJwY08KdKiMvXyQidZ6oQ/9NHRpU1tjVCXYa4axvyoiKsylKSoSBO3ENAMLsu7j+fnTw
tqA7n4wr7OiooblKvsX75ICiHshJFj4u3Aw9q938dbJByuh+6crxL5bCBTgxLGiTwoEGQQ8c4YpX
3tYwDqL7LE9MA1a4s+5Q/RwHo3MzeyWOFxKMCU34Rf8g58+ttRV85+WG3hP1E54jvpLz02jbgIsI
QPRF/908Hn/sX5RVtbGUEjWFVILVfzWuCKxmK0Qp4ELyoRx2SOfq91lUa3r+Bz5nGpbyNhsZNgch
Ya6C34/H67jHg0U3J0hOc4JbvmYhwenHj4CGCNAG3Bf+CszQhsptzQIyEAgMHTX7v+TYk9RRoGhs
o09B4O5ZmbGD3lp57k46Ac0W1cQXPOPfEoMbgFNgLVCCmc3Bmf3j+G1cFkU+kuWIFmnMqllusOew
1eK9OgRPtQc5HeCamAVROPgdVxRy95Occ4YDXpyjD4COdclw7aHDUboATArzzpdv8oHH0PUzvFdz
FTRSYhqtL48KXXJjglGaHpQUgmyIKpVHDJfTLfUokoH9KiytLWe59n9oINq1JUehClE+5nlZ35rp
2qenVMTndP/9hUfXlvJ1rL5A2P9A0icHAs6pf70zlgiCoUxIfYshS/STe+nJ8IhpQgx0/JnnnlNF
PWc31p5aRzeGdQk6AsG8iqpA+p1zfxe+bVm86n2LXCN2hb4bnwbq2UmwaL78oKG+3sy0VPTJJc6Z
I63EVLc7/uowuaOte288NCfHQwYgTTvFB2DkEV9gsva8n3uJk7W3WgNoeJ5URaexrZKJTO7Qiuxh
6tRsgdUh7Sw0C5TvuuAeR3wOQ2rpLLT/xb9RpIAN1hdzgBnYYgc+b4sRdTJZrTMf03DYrjhMvbmD
O0q5qAeAa7ffFVvrG7B8i2Ebl23pPyzELjdIbXbZpYxWTurDQYSVi6p3vHMPbxuIpCWxR7F18h5d
hjRUzMpfeHhS3apQkS3Y22SCuiv4XOq/WV63E8YsBwysgRhJeiNsCtYdzuJhKvg6EZfSBfoHrgso
DDcBRBxlBA2O7+I4IKi/DQ+ZId2gYkkEPBxRcnNhfjDAyrIjw5lMNWxhtODhGMscJwxjl4kkUtaV
fuQ82VsLQSMpxJ6/3mUluU/pKuTAm+uUpBrIw//9J18Hs7OtgTo+xjlLp3tMpyNmwivyg15CQyQ0
0OygV37lQg6wEXNrnUkbse+T0xZolEYPKAwVJVdgTK3HPTyFnEEEvb0+brVpUQxhyAHJyDd1zFDD
YQ9AAK0M+m1zdGkgv5Jv2KdbTkS0D6zWXu2+xCwNm642a9bR/6kuz1o+u5ugiKdpg+xcWSEMR15k
y/rifWaKroUcM5118sd9gyIXUDIRbuIwV+xC8/rkPdeaCiuTFguizywAxPqraZVmxQomLmh41eEq
U9L249FG4tdf+98LxozbfhIcGiIk0H9HrUCWsKrTOeFKf1BgL3dG4PaIV4SMAqp3LIu2MtMNwOJl
YnmJa93Hm7EGTp5fCICXLqFVfwHzVe9E6LbBMC0ji84AQPr75d550gLGpojYlwboA3rKPDXtKy7W
43CNwz6SEUmaJDkugyzMnlXqdXatfqXixE8ANUth3q6tfpt52JoBIMv9K3pCCa0C3++j75pkMOPJ
4ChVDsWmASXSgDQGg76UxV36GK6+t7AJionLq5oxRGWt/7F4BTvfV5DKrX+gsIoJyY2S/K7rGsee
5H+KGL9apXUZPnHFZThCTMqdQYWv0eXXPV1suKV/Q+zgxc35Cw+6zFVvJJfuj1kgQACfLUgOt/iX
HR0bJ1nhr5gHJm97CVq/GMrBfLAVWH5dxjbpjj79RjG5S3b2BgQXmpB0n4yQmeh0acRVGGA41ucb
FGHc5YAO15RGs/yavEb58XWVOKEjK1v1vXrCbJ7IrrFXPBzKXP2rgZ2tD2jPZ8m+ExI1IFkK2yEA
xcKOeA0MhiWa3fAS1yhjmu5kreYq9PF/rMTBEu+Mgb/wdtLnopyNcNgN+zYQvd+mV7cBMnTSarbE
Tdz4T3FwIcIymplxVli6GwIL1tni8U1RJGyJ6BaB8xNVDUhc17+cswk2lKAbVJcX1YR+9EcSLwhd
1h34mqUbOQ5VF5t6wXuD9HOt0avmlXt/cHOZEYZMy8oiear7QXOL5uMWpzLny+1dRDDAY6tQbMiE
I0YAlQovvIWycSCA1WaxesbIji3v0NerfQ0pcWLmVf29V0M/7gULzR9pD3qVyi8he/75rPzpC6pa
Sm6GtSx7KK0eSdbCqUjUQJF9KgMvQej1kkscFz/Y5R9eNuz7JA2HRzg776e92WwOPGye2ns3eXRD
MeXeGaZzTsTvRuqhM7M0yqVpx6vJ7yDziTHj8Y2prMynkBRTGH7l6tFoUZRvWUuUE6gKkz9NPdLJ
odkrTzvBOdBB1Ykb7tYLY8cH7PnNyEKySDOQ3S4cBHvdnz40qNvYBTyEVthM4AUbZ24XwkoVFhHH
tGw3Bmg7Zi0v0iVmG/I/PzriPjhHixHI0mgac+bWfT2WdBw9A6n9xa5emcuzAUat8r6gCD0htxS7
485f412s8M5Ve1PsQPvBACc/D8FnnnCpSr6YrqOC8DyOnDuAOBChdW4TaOZrbIY3NrhFlemi0K+P
aW3VU1hsfEdYUknLXXo//QXdngMjE3uBHma7hoRbPtNzDrb7+jGCAhJBHZZqRXTI0LTMRJCNRKXE
KV0jfpNkaFvisFnebClV9B791vV3wwKDz2b1QQyBFabX9eSXfSzZTA9zwpcnhsPC0aoBcHcXPzYv
obxG1SpeU0mnAyu17y4IHQXkJ7/d6bRfUg3146mysmqJ/fhaGGW3QMJJF7E2Zbghyzhj/dkoNJsr
jK0ZX9kzoiF6ETCAGCTK1+gTNJPPanccXxFbNw0DUfXcNrc/dbgpmg77mtxNTJPWvAnkUX9MOYp1
L2nTr+lXQVcZWOg+E72ndsGNR2K0R71KZEkktxpENJM0j+DXNmgezSyU4VEbH13LTZjCyt9yvclE
fa8wzbObw+aztI3tIuWiqIGTZQMplN9M7J+X9qOtz+BzEqmu2OavP+uD8fM8T1enXCjCMj8dmiIz
fhUK6nB0L6y/TKEojArE23o/fDPjjg5stOgnPMC1iQVkj/MtSw2HxGE01hjvfRCeiHyLB4RoVEZI
s5KJZmcWgAZtRVr4cmS3gdb98/ZGCK6ff5jTA5rLic7cJ0MxODFEtOVJ2EN+aQ6xEzghE8qHGuSx
PbGnGVPGPXnWfwUcZXf9jtC6bPpB32FE9qaPZim0FzYyYR8UX6I2G2bUXBxM6edOA0GEOM7wNdkc
qka3rVb269ErvSDKUFqRlnR9UUD8QoyyDdznvTO5MYYiX5+RJzGVQprHAjOoVbmzQqE4KA8kpQLq
obwNbL9MTk4MOZhiqzcmaXRrHfoHhxr/y4V6CgQA8/VVjBpcato/bLvCKIEqYe8DxU0hGKK75hYi
y4KgOdPuEpi4woRfOu+2y0WM7Rl+07QnrP0k9ft5oQNf8/5XWZoDl9SmOfCBneJMcqTTaSUtVBJ6
CXWIJ4YqZcyKOyEVRvqLfBf1P2PMsWgEz0mT/YjMehS5iViyOTMCJBoBTXb7SylfjVnxf1E41gfh
MmarT6V06xfulSBCnroZ181Vrd9qBKzhj+MJRbgJwDwBMOT5dl54IuzE3oq11TGAarGO69sO5LfM
ULKmJv1Pe3REJ+yGjigaWnlrLMoKYIccVR+Zmm6xU6flJLnMyrKM7F4yb6FtmM46q5xaBp068yn1
vcrueNxAamKCJiSQuJmxeQxiHMnl/gU8LFRdrImUEWY8B7agkTp1BZ1lTgKAMZ3mqonU1k2vLtj0
+dTNCk5Dbx0rMXXpb8CAp1Z+qXVJTlI9rO90gUZb+QD3k9JWQqLq/TO1+jgVLj99UWsxkyfgIBrK
yzzLGm8MGkl1zX3g+Ubq/Ey1HDedQpIZ7ZDPLhVP7+GbTPUPaivcAA/e1Uz/uOLn6sz4lT7lbUal
P7yfpuG8nPFolr6juYob741M9r06h4N+ZAg1EBw54L/4QnWt929J+9AqjBEVQuclL05CRRlTrPli
7VimlAhlwCxrhmD5ezI+9zSrcWCbdxtpM2VssNzAxOxINYDgjljeyMVL1i1MGQu9D8lSmrjWGcZu
xNA1tAvowwUuLUqOkmly653Wk06qjL5WHOiclHudyEk5ixC2uk0L7+hsL73VV1YwSLDi1vgRVRgW
icEqyK23utMygIrZIzcVOUz1GTwR/Qn0j231GJM2Ia4u/Kb9zjvsABZBhBnkd4GMB841VStRJMip
0NHdDbqjyMgGrsBEuiRwaukv/yU0dPjxQ9MisFBAvn8TMdnpixFEVfMezuLiehw4Khw7nWnX+WOk
uq5tJc+QT87F0NiR6fAzZni6P0Cker2vPr2Eg0Y3jzMPPbU9/A3nRrwoE628QaUux2OphbNQqj8B
BDG4etah/zY338EYHQAb4E4XCqmopaHG3CvaXEztk2ZFIL5g7vMicCCw3v0cDcAiTqjlUeu0jo1I
sRkd5bpY2YC3Car3LoZNq0WQpvy1fnzivqG33+lkGyvb9ooSLtbvy79JG7I00JIs9TGWV50Bly31
5R1CVV067UYfx1P/fYW4ezTajywO1XOz9xS6HouIFVMdAGlUyFVQ2kJALWOd6ayjmFZukXfJOepN
c9O0BB9FhRVBRwsb8Dpmx0X0OcqQH46B7t8+Jx+ZDK+cCbSYJeQBThi8U8hzQT/oMMxcl0mQoPA2
hLKKkb6JJmTMP6s5kx/p6A/naluvHqbvM9yhVZgggVZolujiwbpVOkq0/DQRWi/pMoDFKj+0uKRc
1nnsPMvcqxuiQhXxbpPEaW5CKlND6EQ8L0708rTUuHxMWUMvG7sGGSwEKBfDzP7oNwRQZBNzSLuu
0cxyGF5BlsDXJwPd7JNP+qQ0CPiP1j5K+GDaIFZpueEwZiIJeMFc/c+Q72Gw8SPGfsj5TuoQRgq8
krSZkFZQ/2q4mvOCC5p+fHX5sgkSzeYWsArUXwBzd9LWPkuqgdsq3MAW6UZg+P1AuWeL7R70tccU
PTZbKgs5mPK/pacK5Hr9LoRU6n/PSu42O+7FIh1gNrEBzTm8YaPXMWs4m5dKGw7waqc6TExsrd3j
DrFBfdWA0an/p4LMY6QBQz3ThjN2QVDebKPYWpFh83JwEi+rkwReJom2Wi+5279SadMqYHq8Yk+q
FQXrQa84LnZQAOoyc9jY7iz6Bc0ym0F08KP05uRIyBgwj8OAdbWu6QYWSNDxf+hzXXtAxRdwm5Rf
EMwvGLXmLps105XkZSx/xhQHy48Yy8M/9x0RVVJ05cX0D1EhRIEPc9Rvb+EUqjjJM780SqsyVRSE
MisODwiWrvJ6aLONXpIkgV5a7l7rNLXi3XATfZWE1WuPIlvnlYoZfhH9f3OFGeQKzXklSCFZrc9O
ZlUhLUSg0lv/bZwJtYkZ7KaFQ5HYeqCTjuiM4otqIGUeR/l4O7W249ojoj2KMRfCIXkrRdvHIOv4
SqIekamyyFTXlRcXudhjI4030Ynjc8oBGHVjEQX+4oDK3UW1SA0gZf/GqmXyPMTqr43+fZ0otF6P
wkj3vdGzZLXOoPGlLV/AOquLogppxA09aN96Q16G8w7n7jhijbSQ07eYJghqvLHYNT56KEffqZpR
MaCeUDkBa23SXlawUOT9shmFJfx+AFolnSqCf3W5NTcla1CEhxwFiOXgAGGoxzWX8K29IAOIv0b0
FNPXswMQxW+aCz01//ChZYQ1JfXB2wF/yOZ6Fu67Bsd2LJdMuWjK+oLhTzJgbsIDsl6WS5CMVstw
O5YZZUOXRp/PnTM9eWJ7VvLvwJybga/OySnzPX65GYZMzZDQfg1D+ACW/K/xz2PtkIWqIbgZDs+I
wGesYQmUMalags9Dp3khnggQGus4IW6eN7rGNHGF8ts4+iyNvWLihF1F7VySQ7Ebgc8HrhNdXL1q
VVnPO7IpVNDiMUgkRwmWmlYdoEMn973YF2r3HHwfKw7TvUr7sa4Ur9QNkijmY+ug0Tcfql1BI2cf
obMYmzknXT2lXw61Jqc/mKCG6GP7yXMLwL0Inzl8331AKEWGywgyRrnARncczgKv31PD49VFx1Cw
EtPNN3N3mItHqlo2efQnRtIUro92ka3lTfQnhNdGDVhCr9zYR/w9lVuzjkJqSffHsd55QZyYeYPV
JIatn27pkgZ3sO2847nOeeF4+6XOjE61nICxVDLn0D4krUDQIMCwByEAaoJuxagE2vBr8Rxqk9tH
kH7ta8U4tsbVMi+c9Z7kX5DG+04wv6SdfChM2g5TsSf0cMTbElxSBU+Y/EDnA25Fy2oy3ywhrFD5
xigQonwFtvWZ3tp3kd18UndCoj7ukJ88HBCSB13Ecs96ekP3aT02Y52GgKNDdoQ/BkLRHfXLd/8P
vk0q5vpHPzD5VZOmzaXzYXUiB42vXiVWXewgpz65QbeeKCa/CosyOXSKnAWi5z7JVNoNqW6lehNV
371mFPuGk6rC3iYL7l127vRNX+Ml3aMsNKnjWnOhilgNtXtgnMxfB1yWlydElFm7TT6O21wq6Z6Z
uWqjUIA+a7oZvvZS+Ifbws4do6N/YwlbJ6aOyc7lGo+Uvidcc+2caD9bejUQDyE0gzZbhJFx+A+D
1uAf8i+AIHyzutu46B1FzKd4+GnkXN6gD+mxD/L2LHyIigOLcAsCHLwAUx2A3XJYERRSFJYxDJOr
P2gtRIloCgtYNy8qhqzI4qbJWPnZ+B2xlNmAah+HxOoOcqRL7qZpRhsQrHCtwjOsk8skbUNxqwHz
ZfQp9T38xwtLFchK6WeimDmZl0ZhQyctz+vhCzBLaaQgxKDDYkIKVzydrYSst+LjmOGasM1GVUHZ
wz5RprtmrKLhxVRPK7YZcoSV+vO+4dAHGy6VydicIRqOXI63pLgyHQyqefb/cdLhDtfh3XoRhYVf
TVPYpGhlbxONVIN1i3fzdjTc9/6+U4bbgfuaLn8d97sWOaPRPAjTIodRR0DbiYrr9DU48Uhf1lAR
BJwOASuU78mmo3728xv0r5JKSbZJC3AU1/j82DiGltCtvZ4XFZwB0kwwj8ZVlN4dsinTJj96tSN5
YPorSqvpxf5PH7eIWX2U4hQtK9i3aU+a9zFY5Say1nrrDfAyJYhd7Ja/TnJf6JvBUs5Pla2RvRyc
OCMDcMR1Hxai9vlLbUrOxKFAD1i4Hs0vER3oSDBiwr2/c1G9Kj1A07nQk6oampIEwTeTSzel/8Ib
gyKCUt4wHS29bJ03v9LFnSd07MCSnRMhIepPDLST+8ZARojVZv/8f0CZcAs1WRquiw1RdR2Oj4VJ
0AEA+PTd4wHvtytjFjwhS3K8HSUTYDHGsGnaGtOwBNwzAcPxSxPMDFw0EiMeE3ZRgP/k7TWvyyPZ
3pHWU0C84GJ5DcYjWZ2Qzly6tAVBbkLT9Rla1Fly/mYL5oRoCwZAmyAzNOqmtaihnFmrSVzbA414
ElgQFJLqOuxxW7gA2QlPuXKsvcuvSLN2po4R7bw/iAD2ocyu/Bz+R5PQ5vRbyLV8hkA4a69Yrk4u
bmcoGBqfPHPzzUGkFd+q/v3Mj9ikBkbNwJAcbJQO7AzZ2hliipv3GLfxaCCQFEr2MDTlV9zKJ5Zr
oKzi2Ijo0VZSyeiLdi8MnOgAPUObQBrPW7Mlj+dXhTgnWQtJjVj3AOARhBaBqTA3B0dlF7TU6uqN
w3VT4B+YXqJtcXIFVL6pB8l4ETE6kzS6rhNmidKvCEY0kSMh2ca7mW16ZMUUOXVA3gYB4PTRuGuj
WiiG3VH6Jwp8swti79o32t1eXmxRrlSWKY5Kl2wPCINpITzXVSjSYqhKkAEULWv4JiRv+I0XtKc8
HXUxOvISQYCjlRedWbIpKUP9AbBOigr9s78l+0o9Fu/rXuGUc8E0ZJ2x2l3YkPsImGrE3xy+PwTc
7MHGiCNp4I9gygyPaU4WfhiYtyQD8Yn9wUnmsb5xU00+/cDk1A1obVBxmmANpwTJR3o5fMTuJUeX
ilNiN3Cj1U7dLSRw8fttfiLPbB+yfwMKoamL6Qa7vC7iz1+rQESd+GqFMl+TOK5ducaF0USOQo9j
l4Sq2M04JElae4UP8N9cZYZwMPD0RlA1zqqP6DX12+vn7QjWp5PpIZEC866ZEE72ILrBp/9V+7u5
XLTPMObh6q71FSDspk7/YK8WyfDBM9eeNb4BFKxzIslOIRIWDbPxjvJmqHM/HmdmUc3vLm9Bugw8
OroMpiaZphAhZGlZN67iRz0+6Xm132/t4WOBrleq6Rzp0B3O8r7fTrYppDt5pLDPB0YPepR0Gve5
K8xTFv0x2stQEbmjlM6DTWzK6DDChGrkXPjRBNtciZYk0FIhfaY14m3suP+INKsw38tSB2in8kCE
Iu7L03bvnCeSmt7E0OMnZviCP07UmtL1GRqiVljYDxM1yyA4P1NBXapxxwNc1H6tXWQGK5eMIgql
y/Le9x7rN5oc0OgbD/fmAlbXWjxUDrZ0N78ksNvevk1DWYYhaGr6Oz4Qco1wqnY6TT9hcl6YvDZ7
oGPoC8NEMraGALqoNWgoo5skXYar8B4txUm3Wb7jA+r4ItaTRDJ1/FF0qkRVQ3yZ+aTHMfVVC7U/
HK0bLsPRVS/KkGNqfvcB8+UjqAK4jp8OkhSS6c8vKv4G4nVz8/kwNp3PRiycrEE7laVlzYppLF/S
GKpgVdHjpVgVzPgt4P6uwWcS/2qIxCmh3lm9Lp66F5n69hDL6PbtqPHWBXx2PC/HBc5YQUz377Ge
zkEt5S95/Y7Zuxgt9XHCctyAkbLUyy4Uz26rb6SHtlVWDJ+WuBQiNFtGVuDwJllMSPigBieNMSun
Q4CJzCjkhMqWxUXG/CLWnftFXOP8Ao/87ugT94xKcyWvyrURLBbyBkl7X+jO8ijkTysL15U3merM
fMDMgQhSTsAqxqygH1mwmjyFn0JOJXO9dUXcOAC6wGXlSoQkQHpOpQM8OClfz0EJ3pWxJ6KQPux/
XDK3BxIurCa+Ag5xZhWvzEDk1BMKbdvrQN9IW/SySvRiNWYeaRFCVFZvW8hFXYfgBPdpOhvfGW5R
sJHCa84KtHZ9/CNyn7jwoG4k3QTtOptp6lVfCux9txmQodAVWD7mWbdMf9zV2CWyLwR/9MrcW3G4
8JEYC4Oantzmmk+b85z4RI2+BWajjpdMhIjpqcksNs1FODIM9STXiz958+pPj0xZ9wog2Do3CxRc
8uK2VG5g0H8dUG3trQshDgpydLL5r+zJugmlcdBDDwawQ57AYlZmwkCt+jX5e2gqfGrL2t29rrVl
g6XnBaq4lcUcb4vKlskJpd5cnCrdyPloIS33OeTKMkONrZ0/0NwydckVuqdnLQOg+TKo4DZWZfPD
3R0joryOkWpyjb7ZRHOs4QngihfViMqc2zUIP7yeQgj+WaAZrLfA+J1EQNmRRRD4j4mQJyT3y9kU
DIqTfeTDPGzhxdfkxehSGCazwnkwP9LugUlteM8RYSWU/QiLel6MWIBKba2TlDnrlSi+cZbatsbM
QhOIUrC/zCQxtuyS43L1r1k66lJQb2Z2Tsjcd/D49r2XnTbu30KuWfbkdaJSTyngxANMoewKgz/+
1e3+YqqjqKoskGULyWJU3kHxS3buUCwNuS1L4jo2OWo3F+4IGkWvwvIRGagqMmZyqLskliBGy1RM
j+L3x+TBNrJYCaO1LE+XQJu2lwI04c82pQG0alYLd9RIC4rCDgrF3CPJc/BtUUij4DSFxRFUtV7u
TCEwvQfdqra5ztWVKKZ/kQLs0Xp+ZZcZoQ6Ygnc7Nwtv54N8toka8GaXXA2uQhKMuDYehsxlIoV5
nvhPsQXTRPMECP+JyhteBbbUPF3VORPvmPhNKyNTWN30S0wO8DAkQRDARDjSiizrXtZvyzmF1bhN
GURE3/w7opXOOlJoMf3BVqUEAxjwnnnrxsl98eNBwnAufiYRDVOJxr8SJbPh4zZlqnDXrCUvXebS
sYnpzaMVscaCuRXZta5iJYU93jti3gZvhRI+Dxc3JFvAEJY1IsASBZCSjbDtbJJl3jbJyDjP8CBn
QeS4U9FPwhtB8/U7IFtSuE8NGqyt2AOQFkLbYy2UixWzciltZ07GmBhQARH9WmODnANMERRGzao0
GlHjKP04LBeKDnyjzAZnr/rVdezCrC2Q+DPFbxCvZcJySY9LTTbNqmyJm/tN5OqI6NUtwqziiWMM
Mb/WgIEmBv00IdalIwqWJRRgavWH1ZuHIh5qXh/vV2gXDn5buqNlP8py/acx+BghqmVBHhyNJctc
MxMRo3x3P7NiF831nPCmBpulW5BHSG3VAncsWm4vAV15ZyN26FYeoebWlWwJh+p7FsG+E0eWLq4s
6i8ahTxfUU9Ca79zEZz4oAomGIT7JsArk18xrawh0jKkIMpB5knbhfPA5BwwXnBPEBr5Fo8lQW0s
HupYUBXC9MPlgX30Uj/Qt91XFON937Yy30y2Qh18/ECZY8B2JUDU4PIdSsKFlS6jXop0Q0N2HGHf
eCRxZsso/u+R4GbQO3fhz2F4FCfzATTJ1UBY3UL3NdNJHyLxBq3savYUP8LTck3ebRQreEB+36wM
pcGkH6GjMf/CJTAktH1mEor9lB8uXJhsPdRyzeUFsnQ5lM88rj/KXS8peZj4kx2C/XZ9p0hHt5FR
lMaPjilrIuOMRZubnwqJrZa1EFvjFFKeG5JMem5pqHxNIg0QHvog9xFVBSmV3A0LR3pUjqlVNR9J
wNcaWO/e0fE2hSw75LdcYxc0pUfVOKZ3uTHTrAOctQ8NwT3K6erYn5yBbda0TD0IdWosC3wPFp/X
KsH10qJs8HoozVXrZC7UnbNagnQgz/2+cGMlPdd+m2+NTccLA0p0ggWZW/TCOlSCqEK0cM/aFYTl
A+nBg0bQyVC1flhynRe0KEq4XXn94tJMWDIaWBJx/QJSeumF2teafdDPnUnsmfKazcwHLRM3uy0s
zY0JCqVtlYdDNZmx6ATRz4QHAY5lLWyXja9K6Rvq0KXZtuuj8GbHy1jZLYlgiKjaYRoNuNsknmf8
enuMCi4XAPOzz5XRcSBsy1TAVjYinE8wdPncLmJlB44raKJHs6QAnvQU3qTT50eh2hKP9pb9fE57
XuMC3diifteHkgeL8v3kmi+Fd//PqHhuGo46oUW04SxAgGdp4DJ5HvZ9yKXRAOC6RxEmLY4XkW1c
enSFspw7IPPYOF+/rJxIIEBkVbI7wRivxjW/JFeZT5IjofvJ6oIkq9Blf1fqsAVexIpzaktJrLxl
x5FuziVBM3pVPXvZZY2mCd//ieoi0XEApGmlZcG6Tz8sR0Z1qjWe0+tWtAQZbhAm4zCknNjOxrc3
Nn7c30gT9WEdvj20hIRrO0fP7J+QQh5RdFvuRtYH4+OCMSnhVWU3LI36CQq4Mott+iXdpa+aHM62
+YxU6FT7zhvDTSh+pi4RZyOAH4r1RB1gKjdcLbja696E7Mi1CnQ4EfgxhpVX7hjX7EH0uUer3WU+
5Nka7DWwkdgya8SmDnn+T0MkNOerhDSGFWvKC2XoZEQUOjP3p5rqw0RdoYZ0hB5TbRF4NJsOITXm
ndD9g7bzuyf1qsMg7xxyfJ7LeOnUCjqdXKtNPIePEBgLMCVZIf0hzcO15U9hucq4yAQ0X8dczwQl
Ke+9bDB/wIk+bD6m+SjFXqQNOsTIVIBrReLdWotcQfWDNvXSqiTIu+/a+T2UeTUc5TxDT9Lo9R52
slDYU9wEY2bB2244lzzC8XpGsDk/2JgILAwFODpW0a7Kkv+yP0dLcyXTzLJUQqFZjl7X8iFa7GKT
2Jth3OmQBL8gRgdWurww2OX6xT3XTKY4rZkYFn8Er/2ZcFWpEFBo+XDQok4VyunEjfU3DV2FjBGx
zubDs7I883ManwcGIPH1ikTVlEjj4l+jsbFwSamTsmWkrXFFM4knqKCMi8VhL220gironol8XkeG
QwDzY72b6mA6jIoJDc5V1+v5RQ+sQUHjFjg8b1znw4bvgjpiGTRkmImbJkliHEiiy/6Debd7Zuhl
QRIJwmmNhgC1iW0M1LMF2YXvXPsKDpwMblIaYHnExWG/HodtO3zQ79LdXXUaATFKpKO33cB2CXtz
ot+D0HkahS+cgoIKj4J1hgGR8DXywuZnQCvzE+u3rgXYu8qI8KcrZTwb8k2e/4+BDlGYo4A11zn8
q87GyTdF2GIFyz4pVQw9rJU2iWK0ks3Gyb6c/n5gIfppU4aO+2cnMVnvHlqRkeKimQ4lVtd8Rc+/
0DGLlaJxHYb4L4mK0tNK8UjAsbV+buIF4JjH0mHXM0UkelovtTiuWocT1nYwqaWXBbSFMLOkRXjo
0nk+Rtegl1D60Mpai3bCq8XxWLYIAFSG9DIuX5pKS770zXmsvu03/Rl/TVfjOTfbSVm/sgL3wbTa
VNCxoQFWYtZ1NV1yAFwcjM3BSwMb2ak1Lkb7gt7ZljwfbQnr/FFh9up4o/JKdG424uzHdqjJ/g42
DW8Zvyg0ZXwKwmNlwce8s4s8DLlWhRmuLWYyDhhaurG+r5P44DmaP2ap2pZPcoKxAvUV0xCKw43J
uWzR7xpF5G9qjPQLvaiZT/nOxB8xBl45M0hEu/o6CLC9FYbRYYhazI3e/9TM3yms4DkO8+ZhiTVY
BgYUVOCoMUedgHgs+XShJqtreLNouSnLPy8TSKuCSfhUEGRJn072hTSBYAoexsFwphXKm+eHZ9rg
R90kjh5TxYrh3exdTFd9XU+T/ji5N6pAi4poIH8M6ltp7UR75Xxjs2k760E3UpxUi9K1UKRp/LTo
m6J0WcqmgqalFTH/yNmfvfIzRPS56aZPu9TX4mVhR7gaU+6X1PCk+u5T3dhu2Tb7Z7Oi+bE3CDXv
CneP+zi+xoILuJda2fJdMqvaiX0wxn7JxcTDoX7h3hh+QxlUzagd0HMrLB5jWqO8R7sxc8ueIsH6
+PpVXgBWw9GyX3MvA0L+ZE7tFvmv9pfAxgImHm0+kNuF3P17mgzS1XcvOZii6kbNmGbWW+Id3BxL
NzAguTqcHGaxtjVWwo2uT8KPgfY8iiLxpIZgUwz3tc9RHzpYsHZS7tnFgxY95pmm8YDngH2xKT/N
9iK6DQr+5+Oaq5pS5NkAIohG9z9RtdN06dGKreu6rVCffJpt3R/r7aq3L1BLZZ6andY/naMJnLm8
cGTq6Ds52/G7WTbtPHXT8k+SBYXn6eJIg56A7AuBv1Tom3LGWRWGm1eddF/7K11NLa5ELoiJm7Sb
XHypKlPqBhOPhsjYcCp0X4shmsuboQtR44LysMAxVTGZgr/jrzX9C3++X1DqzzwMOAfNMgtcSp82
qB1unm2V3D62YGsq7Id9+mp1aGNKapy9vpvHSj1fOIlE1Lqzz1/2Xv/IY/yazJNrEWfm9ihH5VcK
KWDngkERcSbO4ylEeSXccQMPTYLqJd4/h/T+h14j6bIMJ3OqNRXIGeaV0zHRyoHyBVPs5YxPQ0QT
M8Px31RajnyEW6qEsPbPNn612TLHCJDF5O1XVK7elLF10x/JCAmGNCdqvONmROxMbO9XzJ/567/p
qLqzZisflvE1FecWcX9/DFn9s6k6TwdoDaoA1ZcZ17R4NN/EZHsnSr0o2cO1FQ+MSCvT4LKAYu3h
XgEmhGiGL/btylpNgGWnTs74ImzflpbaGAm+eLeNkZo2VKqU3d+AHAKdFQByJcHY5dZk8MxSlW6y
g7DrNh1YgkBkcXngUF7CRb7rQJkggs0uHUmylUoIwuc/DuHth9V7g/e0r4Adei/TzkMEQKVvn3Is
GSDVyk9DmFqOuhgIq2THxKorMs9CMpeJmUPvtYDxudjexc9vIPxSlM+qneD0NtXthld2pBtk+O8R
Hve08smVpv7vjc8lkI/zSmOnFTzbwgQ0vafTGigTmKh6OGInfIh0XVNHpNiWH8UA9H82XPuO38WC
iOw8EXuFKvQqWHMariBfOYjhljt6pfvvrVDMnUh4aik/Bc8i0NS9O60xs7xlUgeIhsmDaIrsKXVK
rZyvKmYoRENle13hLI4WG8wANpg9FCje5CB6b+4/mZvf0Fz2znbnxHdyeIiW8jLbrhiY+F+LShpz
+1UJ7rE00kg+UI/djapBySefEDQIsK8+ASxT9kwUgUTtQvRcRy63xOE+OvZFTeyHEfucBRWuZ40I
5shVsI0+rs7XGN8Xk7vgpDdN/fN1Ev8NaJo0kJUuq0MFXWdRnT9pLE2b+4hUMPmN1SczDkVH0gqq
VwhURLdJDqPUSG481ZPtZqxXWO0hS/6O4idLR/rSeCjP8fc+O55Z2Kf3zm/YFLYu7bY2piqgCG4W
0VQjuS1BihZ8i21uguylMXpohIz0dPTD0P2yiwqCsaeSTpcXkb2ManICFzORlVAqQb/CUVYzKYdC
6PFpGpru6PDsbO/B7MfEXpZE8+CwFe7d1wvRJOxfJHGFlN0sVaT3u2hv7efoeVIXxXgWBPG3ckEB
qHmtR4/sQGm1CYD321xc4IY0tzcXpLdMy98N1+FwmVYDWY5vFYleXA8Rly3N/qyUbMmep7qfQNiU
CgQa10/b4YRbfaiRBcR9xcGXeCgxKBNTLjGqnjqY+r3Rf6fqCY785X+MjY67ViPLug1tEcH5iFJx
/0TRdHE9Lo8eABN4g7AjCm61GCQGrH4CyrbyKja7BtqXFIU4pgaHm5X70Sy6JaX3kh+rSBmo9NWN
ikm8xVuGQ43IAU3rnBWRN3C/WqpzCM+7efDSrAYfqdHcG8WxgKuI5X8ytR7fjxkgePG2KwZE89M9
NmXZUIiMjkC/UqhDWyRA09FkxGYrMA2AbHnbttjm5EiR/bQWjY7duXKuuz+oE74cYK7P9NsQLlh1
1yv6l9ekIC4dtPP3wBYFbXU8wfpTPJ+lH2G9pgaS2NeOc8iDLXSkeU8/PopzF6c/rh5XrpaSXkIw
tQA7yfSnBu6kHEoOFgsNYL2GDEh038jfYg9F7Y9CXoMENSZ69gD/rWY3cdWPASjG8kWI8d7QVr3Z
iTMNBpl3qM0DyLMblvJV4GXvR56zVl3DGppyFrOn0XrcbhW01sCZOXXqHwNZUPVcGC5R1926+ZUS
HDUBRQ315o8oESMvKD2muWPHbNcmOHN1H6iPG8jYf18gZMxfrGXsiwllKvP+xgpt+sNmSUaHHLfn
qGzFWOAaN1IszAS9M/RQLDfPi1jCVEzqK/YNsqxUywDbRiNZBVcMvsfmhfvNy6E6t2UaOxBAFRH/
vbbV62KQgvl7FkeLvkSUMAHJAE5FdDK174vstEMFg5rujQyVVduV4K76QI9R/u9TwSvjlR9NEy+1
Rjl7sR1jYLDrLtF8ABYGzp2zShCnJm6ntdVzXklpeYZC6R7pmF/q6aMxTRUpjJj91PwzDRyKwfvb
1ZrpxZxvaVuVPd/8f/cIDuaWkh2W4PZzAvgi5ivENogPNFcYTDdZgqSM0zBc8v8dWCVZxmNT+ZB4
VbwEdyC2NL/JLANq0cNYiuJPmkMfXcJYlRGxeVu6rCkABltlDkZZ9BJziCRIdf2c/56PcPV6yTJ6
foT4NzOWbZcn5EiHHLW/RglCjxehee49A2EOsFZy6AKAlxlhFZ9vkde1E2+jnvFB2r3lXF3GJX/h
dmJ13nmnMeUSQzX5TEjU1jycUIMcYvjSiGj6+QTfvvNIRlNOcxV/7rfzDFcSHzcqXyceZa/QkSoQ
5zrmQ821ilDWMgGbpUjP/8QHAhIpWGOaPDHwxRdFqxEiNwftc70JsMAGfvaI4NG6LNqQ7qQv+YpA
mqNqvpAc7J4Y8/mTAFBrcwL3uPmGcUAELnMVgT4fs+BmVkQzVL44Qx+iMNhYoImAAo/yx1+ZlkKz
w+BuyqobHRZOJDw8xc0kY7Vrxm9XIwtXiXV+r7ZTqLmMFx/DnHR6UIaz+2jnLgTwQc+9fo9OEKwc
t019Xvzg7syHtT3JsNQVRV9qgW3vq75ev1IjJkXlwMZWA0bK6cPMvWkGkZwpoBK/5AhNvsPxsmgR
WH3ebLZyF8sxdSJTXfUfzcl9Ht4B439xlXU5he+m1GTIj5mr5Eaj98Vl59YoY+A0bmttU0263Zws
cORpZ5Y6xWrAOwNmUVUjnbpB+mjZa8/eOBRHIXHr/owSTLkIWru8tIcpTRYT07JnhBFnDZ87ZX++
mrW46GvYiaL3FwiBdfyVl5AP4lRunEe2mM8z7zk3uypaS+xFmAROe3nSnhVv/PIEu5rWOpOydwTV
vPv7IT8zNdmD/kRUuTQEwFqzK9wo9Xf79qWe3GANUluEXH4cW1ge1JxSvphvE129oE5fZqe52JPh
XIFAGMzuWPpJva1vqxYJPj69gAfZtPdT9u5A+kQpSDcIIleWBsOgti5PLwD9obAyRfrh061ldYe+
vLwwwFCwB8s6aP4XzwMiLuJMsWeZ2wOunlGGoTqY8WopkvJJuAG6qLr3aleosBc64Yc9wgP150vk
X7RT7PiM/je+MZw35zImdeitPRPqzAm9gZVrWI2nv92mVQiAC0xb4v1buAjCP0dVFKYhAvwWBETK
T+aJTfFM2Te5+xK6tTsfqKIGiRElicT1RVYeW3aDWniI12muTkrTX0kRp+jZxoiYSuGFJu79D5dB
arexYTtkSpow57J0ESOsNQA4bYwRKkv7XwOE1rYSNCAzmAq8kIiDH000gmq+gWQV17n3c1sad5b6
uvGKoTKNY/Y7aSAymGgnOh2k2wxEh7x4mgo0XkksZCuVHUBlEtHlh0oi2D2Vhs2YrtlOVYrOGUgT
cnfirBLQSVbhlJHpgbckRPP3BwB/HHFd4vmAdQe2S/TqNFPLxwh4h+mb2wRt/WdU/p9Ltz1xjCsw
Y1Gv1TWl3GHIq/Y7ba3XWGuMn+woq5wXGfZYazNvOgGJOdqHFXoINv6iJwJTTBnWue0gE3Ye8Xhf
JGWui3JNwCSHZb3eRfhs4CTQbr3TiZvAmw4UpOfgtnisE/R/cBo8N0UWstZObB+57XkWa/ge7taJ
2inxkmY9ZixvNvLVQn58FnwD890m5nW8rvsHg/b4499GFNm4Z+IGsPSQA2MOvAYMImHr/VYJeYAk
VD2HzLxNak200xJwCpYkV+5pMjS3g+Df5nn9l7r/6bEBpSYG+mTuCI8Zf2ZvC6fAh+/vwKPXo6/3
JNOvGLjcj+vXgQm2z8g6fnH2rxuPawewmiqVvvx27McOZBfOMBs0wLDNIBTSei2AzwPXorih03KD
nRdsLFINL1cuuBMHce77VLG/Y9xwpxoqaEax4ZBEbCaP++U/Nu0kHaR/UTB/mojyB2httake0qTc
8oGsZFUcDmOufpQn+lAhNYPwN3c1s5m3Fo18FVLp/P88q8DmEDK7mQJOsUnsIq29ab7Wy83gu1/j
jZ5yQdZGLu/BNL0lmrUpZ4Av5EiG7R17v6JL2Jkpchz63obfcK1tZMIip5tIcxAImciCFP8iiAD+
NJgVGNiJguxRfkxnd133Q2teSlBModqSmtBMr2SH8V6NdeLkXErQmYr77exWczXJlwhI6/yxksh4
kZEM7Op16sx8qSe972H5z/Wxu2k4F/jsSojujHSdmfDaOKCWUmoN6/OQwmX/5ZTAOgfcL5CqhfCp
lQIC7uzzj0sgSVezkdvrcRiwRB8CGC4FuX1ZhdR5przBLgEs/pfOQzjOKhD6SDtDBTrcurSMYU5w
rMQOj+C2b+o9wORVJHWWez3+3AX1m2bdc+/XMYBUB7b+3sjclJWWyWG9yrvTxuhRlCjjvvxNaucK
5d6SkxTiMphfx2SNt0xSxUsv0g+cGfZKa6HRHS+Ea1bVmA8gKo2JdDp0W+c3s7fFGejv9rGwsCFw
B8Mpq3XZja/IOGw4EXPXeRFq+HhWxlsNz/H04l6aBhmCVQZaBEt5+kFfiBj5TYExBB7xyCXduxky
bNZQPh/ucBQ16As6RTOmRX4rpQAcSy+4my2l94F0HNUUda90ez9p9dEC+RtHlovNvNQL3uqlshES
stuI/Olll0VF6En9h5LSNmCbmk/EcuumFZqW2QTour0mVe/4tNy9FoS3CoGwXarMkNuRCJ3nPCKO
HXfriit2y8aBBxEEGs2qbf7MR6HllKD4xbxdArd77or2fyKqsMY38cevDJwak0HOCBWQ06B/nqVV
shKDbnvO1+PXkxU1aMFVsgdxi8DpLBWkQC9R5Wycuw30PbOvUVr+ERq3BzAIxbE3g5Y/Hmr+ihvh
AovrKcZKpQYoFE59cUjCUh4HoiiMe5apurQAVVSI+Pi5o9C5vfxd4qERRBuKcZY5r2bl+UYD/gnw
rOrBvY3MJTG1RBklniEH24yBvUZxKoiPmuU1ihGQ2oaG3O+gdIBpICNpXAb9Y2OTHuospWjx0M8X
9h+j3+HbhQmZKBxQLPZv8cm6FX/3z37yyFM7gHZNK01KZmM8RvrUiKEvWl4NsxS9BAHuqtxjhzTE
ylJRswqMgmoJa4L5S7tk3vffLW6Po0NR6Z2Mpp8SyJIeMqmPz9fR80LD4HKV19t5UQhECznpKaBF
3Pz/0iAlEKQeixKyM0ObSCqgp01C8fC3I/hTUVWC1x+Ewejsx+ujoOyqlpa8DtkZVgaqPDv7mIyF
XuXwdCbNbVMCru59EZ3KGTs14KoJwyiWiYCdknmETFjStoJx1vFm7B2ufkvMw1v2CZSHTJfXdTKs
paN6jPrGJxQB99KU+1cD7q8IP3KmYz3tE43xMjBYblvnBw4kguscGzjrYj/5cew/H6OqZJHReadE
MrFu/1fkCUjmBP9gUHYiQsNZlvadCIDtUL/+hSVYizqNjASL/KC6HPWx/y1P9IP1UdxcvHzl/5PI
Hwgr/F1SOpoa8xNkK6gPlxozhvAbANZcnWfuC6hPJs2REh029k0C/jFgvCyLBNQJECFuswLkh/D2
OzBw6S0m10QrJ1EepIYSHkVOddLqI2iSvHziOgcXQBCm3UWoJFyre0GuSDRro79KztQCR9Mjwxst
tHR5zalCkOk26RpLuP1R+Pjvpp5lA70wh8WG92OSW/VrF+P/CoTNxZNn+YgObfLlZGxYVdULUUck
qUTEexBLufsYpgkNO4+v6Wg+uS1qBc5CIVEEIpJcyhY03piRjhQA/GoAzKNT5OF6Mhr8IRfk88HS
S1xNL9TYfhh0s1uHAiJg8Z6mFaXoVCdKlSmdvvyQNAovgdUU6Z4p20nSIsBregKU5N7ceOGkAttk
TaoqSPmm8+zVGjOyAKynUgMMa4iEQi41L5CzENrccbPp9A0SvuBmM0LgiH6fuEqTt9+wj8zIdDpb
/LvfxT7gNwWC6aJjREtZ7A+kUe9j6aPPkGkQ+m1AIY0q1uqEr3hVPCRlPejPp5Oa2oV8OUEFYQpG
C815AWJeKs4cuntWgeGcMUoQ1L4Hx0c6Eb1oNVtRpo4Js9Rg6vcPKVydYfenpSk1uCRLMKor1hlA
NKNZjuFlppkUKOifMefvobRpIRzHoeAazcF+IJ2wPWExzeutxRdlHAiuKosHLcYynP+WMR7Hkrv2
DwLeVrDdakc+wlJSogQTFQU6inexquVbEQyI/eJTSt7cbUqkVRWwLEYEY9iFiscUBTRRITSiAnP8
4TMQBNohyOHTf5QQUeoTHPjBx/H5y4783pnVC5vzYwUN3iigvad/2xFhQk/+jCoXmPouHWS5Jo3S
sMVHJ5hPpKgi2lWLBeTyKJtS8zx3usRPnH/AK9F2PeQhqiwqAXnjYtTE9BV33Lnmtgl4LzcqsO8i
9x2z9CNeOZjmEKjHO3LRMQG63hr+jtEcXmhOSvd0wU4INb8JFia9LjYsunYVulcoonlmtUt2HJJh
BdopYA56z/p1DAsdCcVFXM0gMQbvesvlYiWZdLh3FR4CKwzs8nNqPoaK/UAmOA5RVsGK8bG/BY1Z
+msOrhF70FD7oQEeadZGrLs8skJkOE+3PCZJ+BfE9Ca4nVPknHBUt6rOW1SeDLH0AV8Epl4X/O/z
GVj8yF1MJftz2995u5x/CWlN1Lh1Cm7dq/ySiO6NfHibRd8gOkVBNyiJl7U0XaSbqdeKhys0jCDo
2Lp3TLl+SCIZMJ8FolSQqKfVbFX5+i73sUF7T9zi1LEa5OmqpHHumX2gUEI7203XYZtCU6aQfHDz
L4FFS4FQsZ96CirowiwM7/M21HBksA10flWDSQPWSXtJJaQaCa/Kx13QAhTTfOzdzoWVfIzOl7pt
O4Wd4taYVg0svDDwEoyOFbeiCFxfYOHvECdTsB+p5yQlC9Mo5PKPx2Hqn3lg9iHrNypeiTRf6oAe
aT0eYzBFWF6pmLDKONFHO+bHL/IPV2YQITFIioyXS7XZe+vYNaYO1lfJnEkjnfvlR85wBT0X3RKL
sodwU+OcjSAxCsqI+o2frngJ0zz2vaH9n7yxFKR71HjiIfQOPOV7xIjoZ6q4PyWx+i7l2ldpejEx
PFdPT+JQutFD8qFxjyZe3y2xNC3jKmaHH5yGDxoPjXBcSx7VSEj+jjWddMSpZ3KVDQmPUjI3peyo
Ae/3wmk5EiwTFpSNCBsNdS5zcpuqgUy66/0NcStGJ9OYid8H+ZKCCu4glTrctoU4CrywV1hbzjDW
6HJzkV63sYgDmI5i8q5s9L6KEOWvkJxtV5WE8MtdX0ZVJA94abDOog1ExspYOBRlwZmrSJuU7vex
XYaedrZfD5qUMjPIUcuIyRByncZSGsHp8IxFc9JI48hhzKxMBaBcVE1QXih3FLneTmK+PfJ0yTmc
Ii2JlliA5tx3mSZL++NqPe1tQRKeY39sUnkwSmkQRVBnDfclAQc4lG0d5XQN6tTyPiJ/CWrkWf2Q
RsgSj7qqKrFo7C5izwG5cID72AkItrVmPbKZyiOEInQ5QOUhbbBa1o2M+cGFIBvVWh5rOagoBGHb
dm18cfcPYpoL2zuAB3kLa5DzERY09GrSjrPpJBLgyzBa48y0NGB04IB5cxtUXywauIsMLLkHsmDR
0Vk1ReyspLa3BHihMPlfHndWyLLDFYTQlyEs2dBOmB7KYXu11ihCm8HC7Nx0pkTdX/jFE/dF55ki
MKfC0mjvyKybwC2+prUjcx6nONkTKDt8wH9qkLSfypbRSVf556ZVV+bEPficDXiExcm67O8rAYkZ
XzXtD1mkgddfwFQXfE2wFbf31F2mAdq5yfi0hFaKtu8oHcI+bGKlNa17LUGbz3XE3/oNjct6Bfjg
0gWQe9O6Ur3TzfV8B+H959vcBthTa5Gv2xC8d13Unj8jVsdzAHngNVw3ZBLVAwWeto9/oFJIjm5e
qCxbRSFDxUdBKkCoxvmmulB8Wb4sR27zHTOnE3JT4BnQropeH5Wq4nVfbvnRMdxACkjpZUDQo+UB
haHESrkQ2kuQhM24Sg5+vmZ9j368DJGYnC/P6PXnYc0sIIY0OzM1gtJ3IPbvbu8X8N0pUoRr6eou
4l/+C2GGcSs+NF0rwLvsWfXRJo9s8L0PB2MNvU5pOErnST6BxvU1xdhzGiaLsX4jETsYN7WUzmft
jTDE7X4tQjfC/o604Bx2g7/0B2qy6XVLscvK0XAooAUcRKosv05JaKYTwZgFnNWacRBMOQ33nsYb
VbqXfwVLuLD4blkAhDfz1+k5lHMmEJsGGmLiuuoQcyzwuouG0FQCUxDFQkLG4BTDdOyrNYrcbemd
XRaaOXNyfF0NirJ1Jp4ADplZEdrWXTWYNn2Cc5UfddGi0gGl4QQ1bWjN8wAwc6lK0atXL6VbcJkS
SZkRLeEUMPNgl/6hBdRnsIe/WKfe1rhpSs4uJJ0nVOBfonMAXL/2JbbGCz5bAl/89XnPS5syv3f2
C+++Ya5MCQw0IeCtNRlDVzIUNfKQkGXE8AXvDyMov6wCw28gaoPn6HfWkKRFIPSMzerE7IhbySvQ
w6eb1buR5vQUvaMnYIj6FWvIxhfSwYglKYZspeGPE7JVXWoYE4jPATTkCtA4jancabp6YJ06mujS
xP2Jz1HR7cO6kSRVw25FyC7575jqkCmWVVaC62C5m+VCPkhYnTU2dIMBI9BlJSa1KPdliJyfpPvH
vQdvpwlgNR1lli7JvSYCGUHXJGvO2TkNpAI4i9POYSNM5sAlaDVFubd02okM7ZKEwHWgY/a/+ICe
WbrnOxIZn1uWyzMusFmsOn3qKnGTMAEUCmWUfVgzwsJ5+8tPTNPwCxw9i0qjiRfmqyxHgX8iS4z2
xROGcEEyorotv2H6ISRz8GZN5rQGr36Ph65EN6F2D8hsxooC5FfMpPJXzbXEFUPu+BtzqSL7xaPb
7MksZMQjlI/M43jWFuQMn/fgExG7EJ1WMj0fb6l2qBG8MK0JdCizQeKd/NpqcGDsls0MDjqctms+
2dL+UIwJvHs93127fqQVacMA2QALwIddeAltsaAOdb1lS0N65Y7ls/tu8VKEolTnFtkvjDvVVuTc
PmMj1GIG51xDUo58JkiCVdjWcziNi5R9PG+/RtAZIF+R1ju25b80/fjFUMD2g4A1W6Xjdjo7OkhH
lBn97em/Ye5aHCGikEXSgOet38BbMdl80V0AQHtcqwXlzn4b1I89m6fC74OxgVZqcM3X0noRfvK9
fDLhe5EfV0/VS3Lb67AgWY0tMaRY2pRl0Y2q140g27ASrobmpI2QKOK+1bf3ZdELys9eVhfVCqi1
V/iRDP8bHN/ZKwJpAoDJPl3lyeJlrdUER+nKrYgWA2hbHMb/cymaWqnLUUPF6egrXBJ9zX3dciiQ
vVWQYzxZQloQ2fzBJtvNTwWN58eWrzjOMTHzDh94LnXTStRFjWfc817lUzzPjZLd323p1CqAdwBp
rqG6aBjkPJmZOXYM4RRQkOd0eCHOuZ+kwOFuHe6Q54VMOBlVI0CVD4/zkLuxLfp3bJG6LTrjuz+K
ir8zAz7SwRXTjEs46lX6oyKg3ZCER7YO9eW87ObM0twyVMiifTPhbk6GwRQ+/uJ9adjlGaHNoMCn
aCPVMClk9DFGl9BWzqOit/RXg7OxujLy1oTguNE0H2gdrr+IFfqadpHvezy/Zcl938l2irfSZotk
2G6pAmWcS700A+jN9mlpgHSzJrYP0KOqgPLYG+VaWOsdKk250HBP106gkM7+IMlCrKzLEAOs9CbF
EKSeS3fzg4RQwfOOfVgkU/QLDXU0Kx48RKYSHjmPI8vptPFkS0Iu7wRY4BlUQhxTmRDRZdhBgo+d
tVlet4k500EwcTsNJBeefQ2/vhsBlb8XfuROAm3qa7Lnn9168rOLxhLul0Ga+m+lSweZbrR5a9qe
S/MZF7dqmAV4/NjKwa7Ksibrn9i2RMIPw2IFHFaZHm/7xemKeI8Isnv+8uGdWK3o7K1D/gVHRxja
V/r0E52vtYrEf9wbspioIUC2JeI1d3QdHKiUDKtw43jssmgwfyVtd0wg7RZXFha88HMB7zXWTyp2
/+dNfRclgrnHsX/5YgIfr5S3x82yutJkm0/2TJXn2uh9R1ir/Fh4p1FYDU69/inKushFQIAkGMWZ
cwym1a2m1Qv7pi6+6DgLATlEO5/WeTWqqpARE9Zxu6mo4H4bsmA9JQYnGFKjEwjYT3+lBEDF/XaB
B7rgBEaGsPc2ajeWb5QLO9uv5LNMQx4782Xe6b8PWpgyOPsNlfyJJrZL5ooiIH8s32XH+WGLQs42
X8FjG6Q6E1m8dT8vI1DJcUOnN38WUalB1MqfVEl3ZQcQqXWoIAUjA8hq7RVDChxgxWfAGZFmqy3/
Mz77gMd+C+eZE2ttdeulFkC0FQXE+CoqM2nGccy+ibqOpNa7mTDCv/wP/QXvXj942xU2jGtYBPxF
4DFBewPgQc4gIzwbwL54YYkPzdWS6Tkd/t40zvN4w29pppArA69QuC0Df12BOC0zdELFr3gvnoBw
wiRj6IZ7yY4M9wpBxMHLT54V+aDfWfNSN4PSHKs4loKbFjURn+1sjnD/Tp9XyUQs4daGjqPj4m/G
lF/m0Y1gjthGAvdG0bIvc35/t+ywl287QUgGuBHpMhMKHsRNW4MXgo48LPI8fhb8tzyHumjkJccH
9V6lwNvgmw4XOXmYySKAzWw3yXUci5ErEAPUvTMvXm+1FA9M3orwkPx2Tq1HeFhNqMnsBbprUOmJ
8mpCxm8ZbgdinKXovmEaFnWgbmc3gor5tlfYektrtKYTngR2+VFTfgwmI8+vNrS7gBH7bg44Kq6r
rRDl2XQKg4EoHI4B8PWAWnqGUJX3A1H+uI0AhHXHxZ7CLyS2qh6ZJrauy2ZZyBVi2wjWad0v9CAo
mvqPVup/PXVAkbymJaJ8bC3TR/WoJFZM8/hWVKmQP4686xAA9J63y35dFK8wmXPIfRsX1H110lDD
oeh4I8qLfggVsfve6sEUvt/+pyEzgRrYI3HdRYPx78TYzMXMgE83YhOB9Li0oz4jh7FUcgbSsode
QE+g+2DQUl+fXTyJFu1js1ngQtbYJWa8AozHWMF8sJzZH8jdi37bYdmuxoCo2ZNJUWikI658NRsy
HpEa5kufPaeEtsjZOfzc4i00VPdy0Ozl50shDjNZcKrrjPsnBoy5aQtb0jrsMGZq5ueCcxYcdK1t
JwVSqCXE76gvsujIHHV9GBnKmKLN9J43w9No3Zz6ABxrGSZBiR5AAyvh0SBwNE1SBHboXL1r1LHD
9mWo2jiKd7cvHpvM4/J0cY6BHVSNzdXisG8kztpvpsD5n4obejllIcbNeDJb+WoMhbfqo2buVwhH
TfrPZ2QdkuHcvggHJYQRPzndFHJ7qOJr63dRo5zChEapz88kZ8kHiZWKfobEC3hTIISU26F3Xwrr
pRKCaNdFF0IGve0pQa2AyuCSA3T65/fY28qJp4XWqbqmc5Uw1MvN9xI/KrTzBXCG2tkt+F7PVFiF
UErXOTbRZ8mfhmLDvoz1HagVaS4SfyaO+KAg4Ea03KF6Lk7GTfbjjYrtYqW2pqftuoVAX6rlnmeN
Y192hIyixISyvvUDbdJ0CazBd6FQd52yjlxeXMvJSs4s8JODHkHwPUqRL8rYdLjq5pCSbNpqM8M8
Lo08TVETWy6zf0jTvhjIbZ8n2TNwL1wONcpUzmGc60UxWzgtzZ/cslzy5zvP1bBybv32hbRNyGY0
DAjk1L8GIFeGxDNHeRAwQy4ZWEcNC9+6yv6fK5SOh9Lu+xDIR2vWMHCXToxdvyYqg4wPe2NLdqiv
AcQL/2KMIWV9csaCygUNLRicuiMYJ3UNdubuFlJF2YBn6oVx5JlmQmyWgmB517cvfiHGI6Z7TIIe
heN+F9rC73ytXSmZesiXiHjPSymTrEuRHEtUmQ0/sZSSXHvmpEP+5MDPUQkTn5BZJwxQCzmJ9tes
HaD+neyB7F2O7U5R6oEy1HpIhnqyANvMiQH6Z0oUIt9tVLdBnZ1TzpxW1L5TCCiTG2WTjL1XWjG9
LMOJNMZaY+JIF6YtUpyUo2ClfULL/T1zpveYOoyIvR0ZOCXkqtDcy4HlYF+p70oaaMsaBwi4k6lh
I2NGsOsoTNUD8/rC0fZyCRTH/iOf9ZEq6UcLZLOnJTrncGVg2zWTA67Bg4KTOhz9RenyO4GU5eFq
mVzE/gP7qLSIorBJNeyam7sZWnL1LOqthnl531LrQBlmF3ZkxPvmoqekx3f/Xkfo6DkHYoD6w4kp
fJhkGAYMH0yHNrtwfirJDjcm8p6zz6/e6PDBZuwxrWVbjymjPnrE+C0B/3Rsfio9LazWbdp8YR2S
/46MbRkxGZBr5HEdJTHSs4+vV0vnLHoEU3x2+7TEXPPchCxe6pM2Epom83URSLxKR4EU3hSUSDR5
5pGvCtG27KDqwenp8yXBDX32fDu4txWz1OpOyFc3kph/5r5ihwayar4MPX84pF1XNNes49JKWOkA
NkOkeyV6cR/MZ8CsM8aE6414S8NrfPnDFaO5sHCjSBwoS69TCH/4iq6EyrlL0RlyU8udqJjZkWDA
tJs/HlEs/GQ9W+V7yUp/Gc05NKG0DTyAt7r09jUX9qXl+leFmotuMeaIXwAFJrbavpRgVhYWpLbB
dW32DY/PW7HLoj9kQ0hoKrUVffMHMZW4i4oEFufcl4sVuMzL4IMee6tbAuUPs2pHF5rLagGpHqHY
qk/XKUSMa+RExt2Mju5xKiJlc/dwTMaTl8icVOleCJZobiD9ux47ZZPRnp/YamM+rIUCpu0NqWEK
M6vnkfyxEbaecPtcOH71FgBiQGme7ggjY9fIto6xCvi8bvAw9TKMF/3OG+ESUr6syXiElubYfaZ7
MAsSyHZVnAapwwfhdQ8SJGXFfLbEZyUemAwFTAea6m1La2MF9hf7+7e8JzFKSyoyEJs25W9qjb2a
hVCwNbEoIlBAfoWXjIPpvbrpL3CTaV46y3VPCf2Yi6lCFNaPNslLKy6cNl/EtJbYrJQLMrAF443R
ynanTA+z7HJoDBunHq+WJnHJXz1udhXdA9ARNyR1uyWLpK/ftpWwIAX7mxLhvdW95lq6Q51/bKao
0elCLO2lEbxuPzNHa2JpeHRYw4kXzst4xMnCxYOhXZ7qka28z4yH4xZ/ao9IkAcO7SocFxqOStoz
TuCptxMZCQ1HgNLc/IyMv+SjEWJ8RmtJWnyju8zlNtJ5WZezAWg2k0bO9AES7jLqJfPghxbd6SGf
T5CEFWDy9XeGz0I8TmPgjRpNHKf4Uqq9J3mIISqm5h6oErZobqQ7dnOA2xfMlkDTwuTkD+My8uIS
C9wZt+Bp7btwm4YA9EUjDTS/JV1V9zqR7MR/4MnG37plKZF132MG7ZpGLoZGY/7nVbtApAY79Rnw
oRfZpMhEYV3rLyjDX2l+afUqlB1MHEbwQ2806uTcX66jQb5r7OJMKV9I5GElm2SKdCyms2sWdPdP
nrLbkolVHQ8Fvuz0k1Q8HR0hzIAICRLqwM+AMALsR5axDys00Ht1ImerElfQxbyr44etDRfPL6qy
hkzh/gNjSB8Flm3srUYDADSpmjRvSNW5fSmT827k4MP/91wvu4iG6Emul901Ms6t9D199wscxGQY
yLQ0d9C1Iej8y1ZlplgA3MJvdrw+05bX2+v+Vc7HI0rhKrFeCUfSW+uGIgBSaf/7aUpklVG6xHRb
VINCiJM0FimiBOEkypIh1NwF4hIwQL87C0FUHd2P+3YkBXDzGJ3qZbgfTwJMJDquyh7vEvPSiDZf
DDVXWZOWWyIeziL09JUU8PfU9ZcDEGLB1BQP7wVve4Uhmgm3jo4Y6Z+AiIBSGvGIY+AGOK7Chjq7
NhpK0Cs9DEgv9brpuEnezDJ0cpNkvleRE+dPbtivWfhH/kIicfQckmO6iAskDq73T8tmxAfVfeA+
gVRp2YeGi38nZ3WE/UQ+QbFg54m/7uSUjstaWWGQHgQnLfHAfiuQDkR5kkzSAKAK9/njDr4X42NY
bR/LyL8XWX/YHmDRBGEz4Hnm2GfDzbt5clrigsRYXM7OSBdISa+dwcxC5B6HMJtSKY8Ns9Ktw5mJ
1x8djPu7L3JA6Gv/OgbgaK0+hslvqJ7D/0kuZhFbFlPPMrbQNkIqjVIckZH+hSfQG7bIyokRoFf0
Chve0U9FOgHMApYHmh8f1yidXxVBkmlkt8T4jD6Nz86g0kLY9Qp+dyc9oO6GLxmKGTFAWK0svn51
CEtHsNxvpGkkekiufXMAAXbcUELrtFyPUefhZlZuX1RuL0yHSwcEkbg4xhwGPw5xjc8R7vsxy4/E
qhBQE6tniK6TX0Wz0SsZz10N86Y2oZVE2uv4CY152gx36x6bgsAjrS+ujZjmR08tGsTpCgfl1ruc
aVJ3g+K55g1kQl2yJWaKIE5N5qA7qNI+uVkluSdwgWq4aTTT6UTLB2uLpEPfUeUqbIZ6IjwjJzWB
PhOI8eeM2AoSkj2+n2jiL88MuustZ85TL4/g7Qp5R9RSRnL4ukf2C60U1lSJyBPykXksW9PSV7zs
a7SkE/9mPIe62wSDU29+TJXq64eJDeN9VlkTQRMhirc5k1S9Trt97izBsOKAch5W1QsU89HfIE8J
oMQyHt8lWIO1qLHjyoB1nYoemOIWvrb0tnL2yHiOTiV7U1OVoXjwngyTrgq8cQtpIHSgYEtR9uCZ
+UeKJFrxl/sFy7Tid54j6+VkN/PTncHKpd7Qzqkrxjnm8Xsx8DwVnmu1zYpiU2Pm9lWQ7+A9GMrN
M76yNv+hWba6BEc1+3Esnh1Vu1KVJam1zTpzvVPKvzLAmlxx7KJ4jz7nWD+6NccfeTLHlJ6ucOYD
oRvA5xi7pXsMyKXIMRJ8rn7wm2IDJ4Rllkx/IVkEiXZsYEIF2IGsJJUCRy3dsOxfoTowNt+VbrAC
euJzMN9RH8qbvk1kZgKWRgkJ2av40vCFtrkRwtyeBrPzz8K98Zdu/qCZ2/8ybiIUJh6JsZ/NBIHY
yzqyRPev0smJfWkv/JAOGhC2YaiGAsCHbTvy8/6N/Lsx0ft2ZHE6jLsFwwuVv4ySRU76vYnhaDyj
QYBiUzvbzdsxp6npYw/KT01gebXY7syWE4u73cM3Z/FyXv9FZj6f3qY6FH5FPkfq0sE7GkXToEfA
QtqawESAbKGEnxnS9TPd3otBC0o4MXOVbs5+5a8i0yUL9o3evl0D2L9nJhyX1Nhn0/Ha5pqD8zBk
u80NsYlfiIVH90qpIDzZygT2tZhs7UaUsrslmyPR2geHod7XRBL0RDrzUKJ6E9El5FfyV4SL4DXm
vSs7MsK7i7B+ATWF7covmYzyWjea9XnOnU0jxaqAt4wzgvktz3yGowpbMWywE3Z3iMrlgQrRqw1X
Db4Dx/GWyEsj1yW9/wbV8YVgYO0u7p3TrRyTK5C47QUICxVuJVyE2GqD/P6IAleacRARkotvcPup
oV+nuSfIdwYsraRnM7j4bUUnQdqqQf/hY3x0P2Oivyg03CvjI3Vp28YYg2N21G5Tf1844IpOj4qm
02jQo5AZuhvNINuvRqsmwATMvcQhWJ6XxClRYzZueUc+YiwtnaHSPiB4qZs1Rm4i1YXGSjhf+FXa
PFWhh91LVEJxHyKj3q6VflJCJWQo5cYd2u+3f0hsYwJjNo80bKMyXUWIfgx2den137LrvZ8E5Hnp
MpjHynFahdE3A1b0PsMxdiAruhA9gIzJaatVD5LI1ZWWUpPZ1TA37/bHr+TGMxlb4yP59+w5jPZ6
Q12K3Q7afKRZRRQCK88mBeWg/4D9NpiQRogaKZjeZyCtXOrnVgHOKW78yOy6c2nlygVBiBFC4jNu
rzWHRWHjSW5mrou2YwJfB/QNR/tXLI6N3W74FsZnO9dT1grpOo8Oey3hyJJE59T2cgc1/skAd6XH
V5Cdc5+7HjA++W9ebAFumiB/M+PyyPGJybmLBDeLpL4Xz85+EyT4ppOkqE5VNq/aWmZBV1K5uo5r
sAO+mjurog+xNggCbL5T/uJ5XcncKAFS8NDGZcczy5zDqdJnr8Kr/s6/+Ml34PjdIiMBBvl/GPck
9sModMD6kc9q07VdPcacwaDnPaCsYfzpfeujM6TJUfQtxU0zZG1567IrunhqbCx6eXvGwMzZhX8D
+Fmj7UALmfgbdnWN6xsDX1G/jmb/lS5E3TgwM1sSKKVsWTpyRCOARrxMDkNi8ZX17vlYzwctD7AE
z3XFcbN+fMyDNSXqp7q5G1KEtCpu45cmBlPSzWp5cKdxRdI6ZMErM/1cgYavb2pkKZO7vcnXdZO9
cS0FVjF/OxOapsCPC46Hr1rhYrQ47OmRgBPcsHCKNFBsjFb0MIiBEUu5i0aUJHyapBzrlA+gh3li
0pDarkoaqO235V+g7V+V8N8vi0wn5IlXhSKCZh5MAFjWo9ylGiBzLxoW7Jf4z/Wj3sBSp3YzGtA9
lRih8+5i5QXF/P6AicgrIXNFYhIgMdIKH8Yh8gRlIKtGbbaa5m7RxD5WwkJRm1cHo4Df0ulAkd8q
w1Ief5s5ZBAyBR7DhHwZOzuVHilPnJSUe9OVq/ct92TLGMLx+vtSfmE+I6jroWfNNqE6HRu3GZX8
fKBb2xfDPFfdQZJo7+CdfhjkbB7i3+IY+nDBkd865e9BzfA0BpDVt0IjCrF9hZ/hhsWa4NHYv/gZ
zfcNFZ+8jPm5yder7yrHmP6tgKf36MZk/OlqycR0SSPl3nqlNhdt9IpP68O2QfPy2ypuUXgxVcGy
sBbZcP8hI+hlRofNonnz3m1+COxjLPLTEcN8e1Pas5EhLYHMHtOYjm/F2aobuX40aPPISaWlkVeV
xDhGsdLDBJTgBnrFxmwZdruYX565A95bWqXi50XCQtQODFHJZG2DCt8MEX3sBaMYAXr4maVyvGQ/
NTm4NOaDdzkLDZhzM/1R9AHJT2mmrYa3jYGW3GVMq2V/UfR7/5oj72Ssgo4XQufDzgiNp691UjzD
DZ1zDjhpuTPCKRXtTncLYwG4ikvtE9e7UNKxSaTL33Z4cxhQ9w6XhHClNsNhi21RP/CUIxQ6Tc3s
fUvjqp1DkL0tGpiMQ7XvbJRobDcvimMk5PaovE0SbL4eRRh1xO4mpEPoJpl8P40DbqOe5cKPp23q
Z4eeNcZpq92gppgiot/5uuyZLzdr/TEJbM4ntN4kIKvOMh7O+mZiZXLVbnHX9SgsNmYlTZX5mgM0
eIy4bqIRZcyYvUuD7dRxOTy/nfbbY4w+oQYZzVRBtGn4yntZztA5OOWvHv+rcWOIgoFQB3ivYjIG
luyUgRrnVkQLtR2IrxWvV78GUp3QZY6LJMKCvvlLbp3wVjIGsY378R/Z1V4HlCsoscRm2qGLLct/
UzNhkmhVOV9p8b90+2jLdU0cpbsP1NfIusgJ87PXAOPBne9/jMlVIdOax4sGdPY+PTErN9qoXamW
NZIB5TB1WL00YY71V0gnDH/f640O4vIWlV3DN7xO4mQ1raMF/hWrfGEXNEg5/J8sFrIA3/hbxA1d
IzKWdFN9a67A9w0KSMoIvtgYkE7/T9aHU+cK4KT/st7VdJtM5EV8wwXLnu2+KNeCw3UBLvGOVqXz
kqLr3fdUqsTLMBau9mEqPnP4xYcqE6dRz9MGU+vH4y1XX1C75tckIPuyEC3l4AY4U/dbPwPuLbDS
S8hv+unELrHYbgqwtG2dNJWwh+KK2vpWP27Qre39pnX1ruUZRS/ItAh3b2of3xYjjBChMIjRIhXO
tgsimqxa/jizykB/f9oawucp8w5FUV5LIcUxTJYhs/Jq29zYszPkElipII+7yWy4pMtjIt/8h+Jp
VgGNLCsjwBmOn9ZqTFTi4fIv/vNNbgT4644QMm96kCEukTQFi0YF/yTjCJt51t23NcKorYZMOTkR
/viT2BtdPMdQdsP7uB0QeFYRuWbM4s3LMQGWAnHhPxiR9TwidcLvOb7lGZvo3gWQBWCefnPaNou2
WkHgRN4KXkXxYLItZbGFv16iYbW6UAB+PjBviRfsbstHuf++oXMLbHrZwxJUcW91IowUIH2FFTmO
3zPUVw41KiTwhNJ8dA2RF2CcggcNFy7wx7q20a/fkCikpydD6qAM/MUyS032gePA0C55abVOultI
VmH2wQw6ewwRyhPvsiNf8JT8wKSm20XcG+IIL3YpC7wjdMeH8K57C9kNGxpaATH1e/ibT06xFJDQ
EHmmZjkUFicQuDYmP8iKkW4pwiUyRVumLOosfeqRLzBFJTAYKSEX4pSSQKNnqt1MC5b4uIJYd46s
2a/e8dbz9996BL4udoRDqaH9ubCENzY4B2s+lEk9oXNLmknKCRhakHn4JjCqm3NuAOD1C2qvfcle
G/ki/CtUY2aMtTiTKUTHoxFdyrconL0jFtax+ieR9A0g8qzEzAPbX1nxWObFrc1FdRANS8OmSZ2V
HDaIs8jitlcAI0wA4Na9W2D51AX5bWMLOUzMWT40pCTYFfx4oGg/BpUSraHckL3s9gTGbZgg814g
8qdHDgxi7NVzIUoJne/ShDMdaVy3GxratHTlPKIO05B7ucUPHrhZGw6M2F0PIZjHtyCr/WAVd3yB
p8qLlDzYRdmYRlvDR9ClVZ6yUZAEi5vPLnowpSRmr/51gxuTjY9bUXMMa+Milz2i62ZNCPL0ghht
XRBoj1lIAftm0VPScktnD1MhuzUD4HtzwCF0cI3y6PFB3Qp6oPTm/BzzxzlZhTFqMqhDx32iRFkZ
Jd4yyjg+WwKyLP87zBxtv1JOToL18pNOKbT3wzJ1Tr03ncnoM6s1cG2V7JgGQZqQdB0Eraf1SaXx
cXezm/gdl3bkSFcZfudo9E+Oc03BKHq3T006uMlXhVC5Lyd7xh6K8DulkfhnXvjQrUC7okQGveTe
zM8CQGrJKBC3hlAcq0EyZd0ke5sq7190nLokw6yuK1ajHvtZLiHWZsPsODn2mD8ecDJ7Dgc65INw
S4skD6SZJ1m1oxGSvwhMLTiQDiQ0ehhSE7EhO7f8Yr7omlR7hXWUWvRuXXC875KwUkNdn+zJY5N1
ZhqSes4WTQvJyeblgaYXhC9K2/thTq7toYERw/nlyBaPXpujK92V6GGr2b8T04rljeqYDA73bA6r
/sKbCBwTvbz/CQ4nZz+ZfW3nCNUqYnEGhomisjmvWduNfQaYZ26XdPc1kqsO1IwRtpsZza3/9O+v
mNYpeGQRDN78xq5q90zDMQXC96P2SnSwqfWjArb4YJ3VKGTDrB+fPs31gQ5xJimI5L1ef6SPHyOa
nhe5zK68+jceHR5QuZtKSuhEO155fWmHTi1jopj+m7TUBm1QZXzK8WnFfb8t2glcVgXhvZD2ORVn
nxo8SQPw08jgwK7g+Gu0x50suRYWs/crJhqja717o/wFjF2l0fERE5qKGc7wPRyVYUXJM+p5EkYY
Hr9gl7JS7UNQpaDq4m81dCQu8AgIYTCmvXvgUqqDa45EsH47yK8xlA8zDF8tQ3tatoIbqcHOwQ3y
fPV4Ru5A0PZebiNQbqT3H5MQF+nOBnk7+Ay/25LrJdgEuD2BnS2gB59M5JGWGR18q5OiGdFhT8Xo
TDLVts+KEfQKjbkU/2pSMiUA3IYXUOuziYhcOY9iv7tOOsliglZ5US9strUjfLXaKJSd7cV/7T+5
SKTsO5RIgsq9hMg6gPgyI3uHjcMUlSR6FGJaTbu3siqZ0AVlX/2/EF6a20YG556d8hN7+vaE3KC3
ECrSkT2KFt3KHEpSO0mcHkOfUd34Q8XQ302ga5Q4NO7xRhLmDyssqnFHymcWYROrzld0PJNSrLrt
SuMbycJtCnormB8ftKreTGU0ebd0STUCFplk1pgfpnEfSiG4PlbPLqEpx5RZ8y+DCX2JYVc/7+ku
adU/w0Eu9LeYhjwN4705VSWyDiE9mERhtySmF201ReUus65D72NtroMcts0B+a7FYFDgX319AC+l
TAIvpq4JAp0ieRvmcYSHPRkwp2ispbhFuVR+h5a2/CHNH0Np6QZfClDeUi2SgDU2GsaF52V4x54b
0jTHk7GGWrr0WuXObM6HrDPgDd/tgGIJOzjzD9uTcN71MG1PEoBD6aJE1aXZHME/tcet+tJ8K5uU
YTNp3jE0HSXgtNuVebC3pIclFxanFDeyYuaQM8bW75+CEyd011Lxpvg6WdzPlQAHu0UEkBGk6aGq
HmlUXLaLJI18dVUKOkmGFM7WRtK05n7sKo+gf9etIMt/QqgpRHivsPs4vH+mxNZG4oRNP6JNVvM0
3j0jd1kWHhAISyIoxOFwJg7WggTPpEQjCOszUTqG9n8N79FtJa0tmTwz9vJ+SPRCSGItJWn2y2Cr
mP10oKq4CXlJILcihL//TrahAyHybP63ozXVpt3yxSrnH25Oza5xSlvMrtErf41mh97SHGNX7dM1
yRDPgMDimHygff7IFwPpc9ys91griHgxPQlBMwQFb7rbYOtDSiMZHFA3DS9PMh9uMdFTCcq6XycO
9A6ZIGrWzC/xUXdBqNEA7JW3KO0Fd5Zsb2bhpYrN5OdmQnC8oF3LVrqtDpE+ZvL1GmtzR2xCsJMq
tLhUD09YHC3qC+h9pkAAdYz/eFNjbrkHDv5nfcFw1hKYGgqMmx8qxwvyRV/G4JhMRDT/pBikTdcA
2Lu7W0hEwrnaeCGLMQLnPPdJw9fjWnrWMjx+aoWZMAZnHmx3vDXgAQQJEMu4FbQvmFmgNGc+AJaW
LMtebtVJbOi/sLBr7uxf4mkh8XaDV57A79fJVVDs9ZGWZE5/on2/tT5IIfRYnJPQICr7mU9KEox5
bq6TrTcaUgwLm721kBtBBiY2+kg2WRfgdfbVo1MLGyaa2quhQz6P9j2lsexQ2xnJN+Sos+Ez302u
edHMkV8NT9WtpPa2lfKNuTibMc2jTp6qYgvsmi9DxpE0AI1SIVbeDejLybUG6brJ7FM4q7TtS+Ig
dhiNvzf1YdbWUP1+lKaXSYNz32tRCw8X4bA/58gqOdi8NvvuSY31kIu+73X0EmO749vH0D95Jdrz
w0ZbDpRf8P07eRbi+40g/poECp0YqsWrKzF04VAbONW+Ztrn91mMO1iS13tQT6gilTR9VaLBHMy7
E6zyCt1zrpyG9CSIjuXTTvbNO+Hr4+b6ueZHFncq5eCavnqF2g7feeXLrxzzmI/bC0uqW4wlQdst
VVdDcQQstnwztVtoToTex5NVYUxNE6qa9aAoHXu5wPCSJxQXfFuJ/u3h9DeQNlT2erU0uHkyR6mA
kLASOZlJ3X3Sz37Ea4naB9IghrwLb2cqmXlWfGljvuoLZ+Fi+qZDBzEO0NSEJqDGlFB9Oudx0RCw
Tp+AoQjPN/LLbJL7chhsDJpUHDxkFOoUgmBHn7iCwNS+NXFgSjWXvFsNTTuPmNyHNaunh+KAOBk6
XRVOBPs+d4R5adbo1HRvMzxdKSirjTtmDdbgp+jvoc8i7i6j8KJol7jeh86JXwnZAlU6qQPHnz0b
HgZ97c4wwmCnJCv1nsGdfudIcfKx40vChkdwMMOXODb63vbxwY6mVcXYdTqsfQe3XZ4Zn9lGVce7
UEPuYgnKlmimRULxRnTl++jPTNMJZKdr2xPdFO2JLRjrUvrkDRTHTKp2H0Jg6V/3ALwnGjSRXgtW
AkthMGD6/GgYJjSDdaXQD6Ar0lFvMnO2+GvYvk3gF8JdIFWktomaMt9pjgN+DgJJbqGfymTorWjG
fbVWihVCScDGkn/HVcXxBbVEEzQeg1HwZE8lTxjMO7/Rch+WCVpxpSFT8cL5jIJVZcRZYEcGROCO
v66E5AowQkEv753lw5zTnEcSKmwuYNPX15sHdbQoEYlC/mZTzQFFGZiGjA6YlHKvbZpJkO5TpwQV
vJmbyUZ2CHBt2xH1fmXkyLo1l8Lk3aZwoV461+nMgCUE5UQ0mL5/WgjpxxM4/eQc14+w2apl3nOf
HYLnoiM+sr4t7IcaF4BDi4Fd3prkZIggl2VGUWR/vCiWRdVG5PCvV2Ql7nQJMMXq1JQfhge1UsHZ
swb+9BWdzu9dW6YFmTq+bsrJpb+D07jfrn1jVKdJInz5jrSbR5ChtUcTMt7nE6P9VNCHjcUkJWXr
18UEDgC00xVRs4pz0bS4+8S6e3GjzwLq8lCs3BokB9nSqSC2XVE13+hth2Tj8VLClUZ6MW1YLajf
EowKq+UASTR37oqmYoIN4Ac3xlkoD0JXQoU7PibmvbRPaHNJoSYdq52tFMs4Oj9HeQgEzyOsELL4
sYNZOIPxT5+fdg38YvDy+7Agz/lfKLWn2SwqiNGDI2bGuscCFYGp0ZKAkDJ9sHtwr9k3eOEubZzF
CUkFAA+ppJtbDGT+GVzdl49VCviGcjGXgOsV8xB6KwtPVP4xprB49gSlV2noSjJSNLxCnAMeSIu4
z7Pf0pivWGvmbkkDtxU71keeDgS3Q2XOA9Tk/QgqiOV5lkvXnlPef8R0P6kiRIaKMbOnws/L2Olg
mIsVT4ydaknCipt0SlD54hkVFjsjQg68MJjfa8elfi353TaEzNMJpCClebmvukQakUKs4utlx9/D
AUKEtprNAoKRjEBpLG1BVBCG7EefN5OA1cAsymCGfADDWJANOF883mXsOX/4uQoGhiIBRobRMDDO
arMCXKcOyLUfPCSXfu/e6kzDKNgSdwyLzALMVAQ2u/BexJOxfFMdWYe64P9EnLbJNbHin3K7ZxA/
Q2/uizlsLzPUfKU/nTo8j0zJspMZF/QeAhp/7lxuOge/Skwk2C/EzoPXb4pQPOkFi1/SLH2CSd/A
WHEVOVpOtBV8I0zFBFwUKuZDctrzog2v7AHGAfOkV/wmLGbBAP+KZvOD5GdmKyKktog6kkFnRBbI
+DMyUTzGzq90chpYN+84Pfbb5c9YuBTuPlS84FecoSiKjz8qSGzQcKhUl8SNTHB9p/iV1o6KYyyE
kehUqMjlF+q4cUIZMBKyXnjFv7N+QlJUFQNnJnFlTe5GH4Ag5+H8fA+60yrE7A+IR2qCuU/arm88
ws79udJIzxXZmRvEZWIaXdJbKfuoQCrWOpUcOQawoPTKDsO6EM66MmXJJaNMH8m7win9xRU04bV+
ynh9IAI1wi8DR9eZvoOKfw9j35OJVBBqJfOwi/xd2PX7y9zjVKqPpc7lkDON9myNt+1Tw394Io7w
yhIx0xygW9wc8TanBYrghd2FEV6mrm07S2VzN7wTCTmZ7lGwQ7bIe8JgLB5bSTiDiBZpQKtEjkHp
wC2Q7MqHJ3rt9JJETMUBE/a0I6JFqKZ2Qovy3QsGv91X9hdfWkBzj9l5RIyoH8VdZHOAzOq4wpfe
5T8JTHKq091BNgRMmrNf/VInpgounwKbokHAMd08AAEedruAC29B8SaFFHk307gr2uwQjugEXkbr
F7nCih6HlGktvpr3QUPI/j4TlRoczguYYmpmHjOiLrwejrPF7TRN5cApQsWx+xGGlevIANuiiabI
Xp5IT979UrZvLHRsWizAn5rMnTkcvzmWUeoQtOVmbh41miC3h9ukHEreyfLNvy9V44zRwhZK5fw9
SnSh9oYHuui+zH1MbQKVyqmkpMqJFhPI2zTRFWpnWgTcQrdC1TD+ZXJPvWZd1rdD/1/HQ4BLYhNv
RdUM4+i67z4jpqck++jKmJcmrUa+jSB0Vk4VkS5basUeS6Uviul8kEftavbhIbZToRaUgVKl/QES
acHatIxWMr+wTKJOv41oDKT8cum71rtxjcxvLgVYbvN0BdfJXQaskZalnKiJBGoAGKzE9X97UP1n
xCMa8ifKiV7K5TlJBp8tXKfMiVQlFut5JL0M7SyuEW73x/WXNiSRtrfdTiMbh5qX3GLFTuntQBKe
naxxbZM1W/TSfymw8S8IUxJFcHfhmNmJXB/NdZkUWO4vrK1EoVQgbLm3KEbLBnuXnQJnF6YYHRbg
5HdaR0St8dVJBQ/WRKBX/CK6SgxmC8vpyuejFqaKRMikfJ4ara3ifWXng55YbhhOPT3CfIycmLaK
V5F3HENjbjbO3aWHsU+suV0+ciwnx2MHegGFuTQgIN5BAdl3tU6SDXldCPQEToZy3DwVdlSdCndi
Ke3WIy9uk4i4uWU5U+06y6qcoQPvtWEtrQfpxmc9Pn8NciPQer0YyVdAQUH0/lsjIfTwsPWNqBP7
IPIJZBXRWXpLmb6Rzj8kOFiUvB0HLxasdiCoHGawCUe8H7o3ajpD7JVZJ3bHKyFx80ocf01jHvt3
cYdZcdRsInbGZDiHqxn/VbvzF9TAxnp1GZUVOT2OjpieDENzqM+lpQ8APfWr4j27ZVQuEH6kdq3i
ZFDp/7Y5BLPTfJTz2Ge2swhNbPwKSXOR7GT7iNYMgA2lYnoRyqPrTkTozqD6KoSuth/XGDE3kwJQ
ETywmKMziQMM8VD8Wg2k1g35ND7HGt0zUA+B1holc7nIwy6Ei8FDU6wxVv7OLbkTevPuKubfKj/o
FnlbqEm6NdX44eg3UaGo1L9P2168Wm7r2bA2W/N0hHZ8xcQtRzDbfCUKwVDlvGLDXk5nDFz8EyH8
imP6G2F/fgtf8dIFLgCEPst2Hpk8Pxej0FpfcsISlCqDtCsaqya/m8LRTvOGbmBk+3CNlv2VfJAU
fsXLnKW6lyIuFIhoU7CQHKrIh6FnzVv6i3nPCIJIpEJXbZOA1it0YsQdTUPfXB+IhzNIzXopu7Z0
Q/AxJPwjyNQ3F25nNTZ9nBOBLU1F5pYBNTAC9UGA7WX5MGJoEvdCl3iSu7wiZVOSBo8daAUrCKz6
tvJrxB/jiqh1DPGT71rUBaa95f1a65vxrlsu7J5/BtjAz6zy5RCycF9Bq9ob6y2D4/3HMoDiu1VH
IQ7Rkggc7Xds3aYBAesOxp2kXu3B+37T8kErRYV5RTfTVRREsSJufSWgteDXgq0deiW6Sv9R/VvN
ByPFXuEQ0zcGfpambeIeOTfmuvf6Z1ZpG7L3ZxO0zqYPclCoPlU8V/LbgN7axucKechuQLXv79T3
uKFJV9l+LaJCcj5KZG2L3uo5RFcP8VSw5KkDAgQ+CEdk1Jq1z4iGlonhIsrK5p/K1DH/7nkilc4w
IfiFGDeSYA4Orv3S4p4+9CxJKkDI+ozjGg0pzNx6F09KnnebtDrXqetpBVOmnL1/6WWiqrEnDNAm
tCrYDCQYEf33DjW+c75tTqC7G0Pm3Ec/3GJ5QRvE7BHWWz3Z3AaKOzsXQ3y4wMHsqC2P9V1+oJ8J
ra1X18nPFicXtmbJ+ZEtEIX57k9ynWyvdEIVvsDMYQ3VQ3I9QKOvXjtlCRhVEPpCEn/G9PRym3uC
pEsMa+QYXzw8Z2Kq8mKC1OniCbfmU7//g9izf+e51GnrasBZvwgOMc/xcv2QZ6vUFdcVnr40pR4q
VGXau+BGQrW0zIY/LUwSi2tx3vDz9+dNAImi4VL8i3+/sAsLOG7VfSyNrqwqSOC6SfIftPmW2gYP
VcmLpp6eVddSpMBXUL3y/k105rYTZynf33y43CzYBoitdbKoN7lz6PgojZbmlVzRHA6oIhJ49V4C
EjK6imdiTWwSJN5EBcKJVEyZAv4NpD/b2CoVIu1B3s7ygDBR0Ww/0Vp9ek7bt3Fkh5CW25N7GcUO
MKtBiAy9D1tgleAdTcK95N/qsp8rlHTR3Qw81UES5v3/ZW1/WQnR6/Dv7LoaILY/gp33OukbK5XG
9c4dAYKKvMhmBN9rO1a+/QdkyJVLYBM2HN8xhBfSAK15CO2EOl6EPKCWe5RP/PV1nbq81tbNjwxu
LPzu/4wZWqhiKkvaPjjhP66XCOj945jLP6WOeMFbnSnxqmJ1BDMWKqyf2nYM5WicQ2D+nPJnyjLl
4t4s+pAmCQryXxZ/KLuNaggv9hBJNix0wQ6TtLqebUBCSowS8xb6Z2SaXsCY/iE4F3V4mP1T7cbz
yJBJw0EVaaLTUGZ98jUkRiOFkhK2WNIcCO/+xG824NMBkv3DcNMiRnEqhhsc0JJ/6BZHfEDMeKdt
tLhSZbG07zobu8c6wmgisJcZu7lvWvOjr83m3nzn7gpXN5tUT9q/zpVa+fG7ju3BZgXVF6XQyyT8
qRcXt5lsXpzbFR4X+iY5juPZEy6I/M/j8BcmZVsvSV+tZMevzzfw/1fDFV+IUkriLktEdMOumIXd
IoUpjlSZ0h+LDHWzXIVJefb9Tu6Evd7TN25dfhTMMf+i+a4/n3FlffSzVFmSsKIbl0iWY72fEWAm
MssJ1dBJw6bb9WkzAlBLBwLvcY08yj6brwteeIjxuFvHdZCdnEyh8lnagy1p4I7tNjLMYIp8UUT0
ziZQQ5p06WPHgduFCBX7HO2abbtRaaZ74sx69wXkPpuST+ug4vRniqdfNyCyyJZO4QfCxztYwRLP
QN68BE5wTuZ0Dlpr3hFsu3sIpyaQL6wgU2c4ocNjuqfjA41KbIGzb1FuT3aRzN/7+RBuzHrjF6QZ
4vaE/TK9E2KbL017kn04W5zqyojt05HNlEcn9a73DVlaKWCq5M4dWt4OxyNaxM8OwFBUNfgNVme1
K39fbVtk0DNPXVdT9x+yIZfPYBFGWYiPU9o5w+pnix5TsgXn2kOoDav7Rd+Rz8okREQBNNVKZT8x
hBtAjIR1xiGj9rL/t7EoQXxW+arVJHY7K+OUDgeTUo4u3ywhB5DvBsb97vV4HGpQ/CnW0T1pCDpq
4j1xINvcTVai0js4wtX/14OTmypyVzxmws63lL1B+I4xs6ylIxIt5Q02/60gcddptivxJTgOobc2
doj9bMhp+3eJ9tmBxpsOUi4vpDfWczXM1+BbaBYwR3oAQiJf0zUDbP4VNjszb1z1IuDlaF3dMso/
Ye9W30BaY19NhBImfBRXF0AWh1sESXLMyqaA/k9pQedBO+yQSJyhXeatEp3vEHuEPDCAzx7znQf1
6A5vl04UIk8rejVK1/78xfNRTbeOMpO5sVRNwakMqq4lCtSKKbqNmOmzurXwvz32qw0K3jjnQ0JA
hA7xK+fNyKHB/8jnFMehoRPu1HKHPwyoH/UqxfH0IJojeUnGN7vBfuxpJk+715t0G+bCiSxP8ymr
YvCyB344zqBXrq7N2370SU1OfJcdMExng72IrLc6Xuo5WdLV/ougYMxMazfhRjcdKq1c/HgSIcU3
c9GoURoIyAGcR5rOlILJ+T4H5r/Lp+TByyI/Iruy3L0BRjwwyjq/HrDexH7fWtWH8bBVzlhfJ9rV
GDipRb7EkUF63J6OIYkwJmWuHmvSj/CcWMvxuzuDJobvaxJEKa4us1XhFOD2nXdy5SyrKkLoeLhV
ngMZlyuWWrm/IZE1Rp4pElgwkctGUdnALIhv1XOFD4maJiU6ggsX6betWDCqjN/l3bqG09bizpD4
vOR3bF/nZ0W/8znFJJ+6++4FHKXTE2ZRK6fdd6U8ccUmtc8V3g9J7P/qYPQFeMwrNm+sTo/IBqwq
M50jzgJGh7PamQquXUVYOzdLfpFFmfmUbRYSajuZ/0ZaYvnwWtarNNpqlhdw4POPkOMegGS8S79Q
CqkmGKGpF5eAY75jmHbqPe/DWSfHzrPCOkIuclL6fc7mO0R5D++YeGwghEBkF2aiEpRGBoQFU9Nu
s1nHxxxv99TOfZNs24XUvZOapwvG3v414kKSB2sJvkdgBm2URdY32eUI4X9AbGWcESWcCVX9KffO
e+P5mJwDkk+h0CgDyFLZKm5ADCqBQxV4s69mKd5oLIfOGyPbEfDSwuLYc5iMEJu30s1SMAIcO+NE
aMaisCOOu9PYxyZI1HKg8OYg7tdP8BDqjFNnS79RUspGOi1CCzrVLczferFXSz4zFkni/HQqzcyp
xy8PeGTJkTSYdWCm4djG7mqMVmrAbAccDHABhO9WHRO25NYSxcTxvt/ZZKHV8GjIt5+wSuSHz2J4
Fj58PZWy+DlvHSqtuDWL0q5HwGtsXShQGUy5R8tbHK19blFfMzT9lEUMmO2dhOkNzlvaRXYEO3Ay
oYlojsxLdg70eMhIo/b7lfk2N18oCkMgeTNs5woEhQJ8/dNKpdx6AIbj+PMH99kie1JDMP4aukKZ
eiiGGheeNZQH8T4Lja7cW4a9OcHTk7Gl06V5HCNlN8rY+BhgspcXBsbozktl1Zr9W1r76ezoawc3
Cudxy1x9kdac29CqOFlgqVGpQdrdb9PwSyo+roUbTOQWocv8nHSlBItQmadGr8Ox3rdC/fSVjSfS
Ixq9U/LiaKnxNr2qgqOMPubPK5HGRjPoyyseviaEp8IwJMNb1ahEL7MBPS9HKenVkNaLUjYfw0tB
uekcgh0A6PZ4VGM5PYUy03bES3WWyGEgEvzuIwdIepz2fgGraibZMlXe/V1QyDZ/4MTTi4xHlQq/
tn2unQBVAQNua+ipd1OAdcolq2NPC4IE/Ik2iuQ+nASIhyNXP4DFrRNmwPBF3+YwJSEBpw4/j2An
/7xwrmf/GomVIvo+KGZxw6XvXTTtZWbU2v3jJdcLwZtZ0k0sIpRq+cNimBQRoV1bHC/REpnV65Z2
YXFc/kSjPQst4GkPEy5NX5KfdXhHGqT2AG3GwpdMgNyxRZWzpoXqvZAC3jsOIRn63quQdUAdzDRk
n0hQjxhF0JqKQjiyaqGoP5IfLBaL2RYi+k0uAoNCVBjfsQgN5ZOPPWS9wwt15pT7upmnPZ+VBZ53
Veh7pZTxGrQ/NNkBae7uJ6WjiPIqn3G/WkwqeSiqcaVsZdpjoee31czsZDet7nWw41W9lb6jHkzq
8w4+cDsgDfJpfBnU54F6vMaCm7/o36ksrVdlSDcQ9HuplRWUdxCcqJdWt8j9iD++TkrhdF0AVkkq
sBh5STcNAVeiFxCVErD493/neCuE/oWhUY5vXnn3wnl82dRHXV/phN2mCemQ2v7Gyeyl0o2YJTbE
AJJw1unEJrl1BlRDfComWAt6SHTNy5eoPMVVokQ7i7gT9DvWAK8+qRq6jKF1T/ZrChncVTJAgcXQ
9V3K4/IImERtOqf/H0TzFKwp7D2LuGMddNqJXznFxfn6Ji1INAUY1aPsb5HGDjSb0OLMpIFtJj9e
ShkkXaQ8paCzNzM3tPF+1FmP7HeX7mqQOq0o7k2g6RGRlFtSvvSdzRE+I6C1zeQhJRIJymspN6Ka
OQftS2IeWEcFfnsoYssGX/xQ3g8ELq1s52VdfHdmrM5MPloUN8ik0hsHpbZWKnZx8uhavHpFGxRu
LdP5dKBg6o5FGL3jRCrLNyREiwo4y8J5UeR4eyR1N3scF2w801G3/2bvHEEjLeJElIXimmnUVF+n
I3hAk5lb5X1UwWcV/TO/EhBPZSItXPFbnCqvfZXrT52/h009sa+1h7vb9CneANsdwqPIpXtUEdMQ
NF9YKGQUONi76FXdyhogSGbcinNDt8X1fUsjJO8LWmFnX+u+EG9BbgFo/owm7QKZZG+SC0DEzZ79
G1gVd600Qwim2PO0K5/u0Xlmv76a7osVkuhwkwAgKALTi9lT8g8Jn/kPtfbrHP6xXYoXl/Jso3rM
oVtmvAyVSzciHb8eR9VNnknbK7ZA5N9O9MFp6MRJPaShX2NQxngMu7EyxNAB3zrn3JN14xOWQmKt
yOuj72Cy+0uSn1V2BoGHoS6tihbGqJtzeE3sZA4qv/F7XaeumPoME0cvh6BxZ41bExXRN49hOQ37
FpEzSFFgnE9qzusCPqB2a9lNL1eWQzJVx9bRj7pXUK23JayBFlsyZMJcxI1p4jo2kt0YhWAUjyc4
RG6m1fTG1BSVNvGrdRtStm9k0Pe+VRjWf5YYzmMsIcEGofSw9XqGjODXLZwo9HjGZAv9GXdmgmEb
6s1nLhSh/n40apHSDZ34vLgE+WJo6LO1dl2gXb//0svAzk/4k5JlpyTzJayETHukTzTIcvhwz2Ni
Cv4oichaicGqEDz4xX009GYsb7c+bQ5M0Y98QQZW2FzCsIk8WmdZa/y8e6hNRguXUSiXakx2KkfE
0fvDpV6Cy5w2sJZQOXmA8glPnN4BMywwEnYEXCD+ajam3vP9taaqlZkJPO3e0XKVly1Lx34hds6E
69E00ZsGDvbYnM9GiK1fhyPhbRWcWVEENQ7kBJd74iZgG93FQrIfqtwpLVhi2RgaHAQCcKZy0Qe3
xHIdQG7H8nTN8sqAZp7Hx/8j5xUmkYWzLH8KH8AcmkVifrwReXwlfw18oupOn9FU4HBEo6+4AOd4
P4q04kTWC5pxpRQW70PkrvKY6EWmnv/WeGfXNN+7ROiXL3wR7kZ7xxawfYNuGw0VyzQ9WUPSLGc4
wFd5yvRJw9LbjUFZvCtjUbY1tlEJJqSx/y9W40yfL8rGZhUAq08sIfGXFc2ULr9aG315s7OvuWp/
OFKQuzvffFWbddph/M1+FJJGkTe6C3Di5nePMOZHo0+qWwN0efSfTnFf6fOY6F8FlXdbv7Vtwt0l
GGRqgui2DK1VSdD3kG6u58dpLoSfidx9Lw1ktyY22PcdFmI6km1oUb4JsKmOW8BJvvjOZmfH2SRi
lFFMEA5Enpgbgdh3X8uFtq9Cxb6vfHvSjiXd36qd82uLpcq6iRguTl4orhCexEpwxYiYlGxYk0SW
/Xjae7bR+2xJO9+f1QFLFvFew+SNBEhszMSrB7oACpZ8jfh2Y4aRG5pkPWq20oV+tg4jP93EzrTl
LWGgTYh9CcRhJR+bGHP6i/0FyPnhgXyNIK72zAGdv3dyJF1tNcszfcgozZBZIpW+VyVn94ssAOZ6
4++/3Oto3ESCpnS5brLX1QqLM6Yxf+mfPzMgTu2J0ed6oXJLnzg4wy3uiICdackYg1vLf/TqYKNt
8h3q4DG7IKGCzSdeO4c9BF6QAs7Z6KSypWqhJrR2yrNU7rQzuya95F4bmWoiRG0/XMr3Npm05lfP
U87VQ7eUJOPeokKtn++VfNXxXm9iMYZNCH0gd6gD9nzi5EzQPFclBkBdhJKlHCKs68/tvHaiXt5b
eyCMFEyT1OJZ/rgU7ixhfmuXkqunKLr7TnwU/qfvJXbaiRWcpv/F7d+7OYVSpw4uJXma9lV3aPoN
m13ucGwJWJg81MLzBuDt4xqBliHANhxBu3mzq4XohkVO1kg5yyXyhrw/enQoZk+xsHVknlglfuIy
s+U2d07CVxJJnSc86ZhbMOEJHRSFi3fMCbPwQAYti2pIuFdIRvuYmqU3CnnmoZNfBkCe/398761l
PolW0kaIuNw8JDQA4QD677SkrSULPNokbfdtGDxYGS7T1B4jGKVBHEt6Uv5jFR++XESgLRMelF0t
du4+j1Plk0/vckXxaam1BWIoTu+pv7paSfw31c9VC/cHi18pN2w/+TQIPqdnpRxJ7Ee0jvcisXc+
htBrB1ZYcV7vkxlCggr6BZmMUPtLP1LwJ+Xz9fqOeVUyppAbXMyoSfSF9woThfKFxyUQAfD8hGWr
B/ykhOgE1E2y2y62HuiJFCx2xeWYgIraSrXJLhfHPKrevO0/QqSl/225mCjbfOnMiBNJUpXJryuF
HHDwBXSfQaQ7UOa17ePWHfqVT+w1to7Isi/Fm7g+PSS/uaROZWkjsB9WqRRXjWsFgBKyqDRTcDMq
WI+wExhGL2eTUmSEC2cedecYZpUL4dhHi8CRcyHT65t2LzHm3vhV+VjwddC36zxWeNPtQ2++5cP0
7PpJg4e7a0XZHK56qCiDMR9Axy1ZsqAvuwBPk7wAgiPx346C7Xv+1HzIZO3LcVpkMgDbusYxZuSz
dm7EC0cPP+aR4e01GAVtdC1PtauRtFJ2NzetF0J3+pKoEdhjmALPmcywzBCtSLT6G2bc2E3/CLWV
F6QQmforSLtOOd29w7uLU5+TOnmYJEIMtp1z+98GdriN94S3sFVQayQN0aXE2+8dzQyV3TdhC4NZ
JuMEqUOvhWe6L3MZUogL9abpU5niaTCXLBI/wwMzi4psx1Pex0zkY6UgX7cnjQtswM1y5urOgy0G
m3DoBkp0q8FVuZ7XAx60I6bC35ZHFNFnLPYhoQQ2O2/6RP2+mS2pq+Xmy14SZvL3+8//2Uap5kwY
Hx5jefE39sWOjN2CZTCpXnajyOrQGNR6YTfmIBKghM2Rv3nF76eT367+1j3JfmwXBFx1JBXd3GcZ
UaN2VlDw+9+xEaSZOHGG3FYHHHlXlrCbJG+MiWcq6AqPg3bxJm8pcqxTqIbR8qIBW9UhivRA9PWc
Vu+MABH4TIx/kNBRI6HwnobYLhkyFfQIa5DWwqTHAkb5ih49qkXfTHX0fl3GQMZHI33VJmjOX5+4
O/MYogNaRzYpNw4IL+rR1jawIHrECP+8cZx7xxmPJU3Q3LRR78arbU//DuhT7v/vNr9ZhUy5scRt
2E6OPwwHlX1mE2vtOFci518z69AsKr00pvWwqfcswkQz9IKhgg7OxqfkY9u9Bc5yOBw+/02ILyxa
ONHxqtFwQgTQwf7bJPX3zZzuF9pjCMOb47Sz8+F0jk4ZCODMO/Y7hSfLdLKSQJmz/trIbcS1LaPp
9FeiIIuRC5RF2pYU7O/5o2S86CCyaJhWcapoGFu3f/hQfxrCvSJR6pqz2uUPLyWEI5RQ3SiVBekS
Drx55PL88mdIKaL90V8KwZmMMYh+h4C00bxuV5dYVkEXhULqvtnoSPxolytRuKz5IPkshb/vi31M
R4nGI51US1NPYO6ygC9OKfwINjF9uUBbO/xY01SCjIdWcN14Z5fZHZqesUQqL3DrlJENZ4SR2JZv
pkWU6lf88+6HIIcPSeFLIXfgpAl+5ZPeX6b2QzgagXzWVm7pJNkjNgMdRKHmJ5yATXGy3gfrxey2
7sgIkE7ZaJJBm2QS6BYFL8D2HrT/i3riDS1kDnCMFjfXUoRn1YjYoEcaUchK7i0quwLA8D148Eb/
yQykzHcJE6P0Fv5Y7ENPtcudZnStzL8jeGuBULtCS6S/alrgoMhJk+NYHNOs0oEdMq66CXJIDeGh
Ik/jwGWQww2vbDnHuPQaJSPW4fNrJJma6gB/DrjUlQfROT+b//Ta2RmG4pqufcABWp3CQ8eFU4+D
3+IHAmc7eTfb1pC5OLxHiRPQ4UQefs7Ngqyz0TIFo62LRcpHTm9WUoDqxi4p8SCizpNCDM5R6rJk
FnwtaHVeuAxA2Sj0oKPyD7gJwL8ypDy5NFktW1B6Ekz4j73KBtlZj9A93Y4npWfWyMJforIMt8AF
SaDcYc5EfbrQGGkfWQ/TC7IEvYHIuHp+vqJfoR8Rv/9hH2bskc5eQ8ENpuMBLFvvL4FZDJz5o5Kd
hiH43vnsBhZsmlZrcIQIlKwnd5umZmhqHKtcJDC28Dqo/6tIblIVvySdjiXu4NkquXMnBrXe8VIA
Ffokd9/MKdeBoAERP2YTJnZfaSr+MDpm6w2pJv39tBroUbM2ZXyMw3uy/5W7LFKTMqEvA0DDy11g
pDMOjTcPSKGp2RPKFWUXWE4F1ad5oGtxQlR4C+PNTSbCdtDOf3zVJjZIDscUbyvWSiyeN79EyWvV
FcgrV+PAl+bn2ZCQEBImA3CxeW65JVPouiCWRaDAP7aag9eQNjVJZdoVCnEhJqCCRlr/kMtlMsKU
CSxKDYtb1bQaGFega9PhFp4dYbYpWs56AATrhSMtODuTjk+J8TNYMQTNy40hazG4lSO+23yUt4ng
iYEWYxOp0QFVlgnWN9hJBKilJMbM0XYo0XuytXBn23r6A6MDQBuGTIfyOBibOBvz+i3gx15GU08R
lJddLtcxNEVlBr96MChQm6YkY9+QVT/DQE+SDbtX4h8j0q4jeVf/NIrio57vHxUa1OlqrVkZ6zmT
eRHtvHA616p8+W0UPL5cW8G+9uKxll+z3Brv4ynwADNVZJjkZa/aBwjEWs4b4GpdfYa0sWqYFQJy
GCVBtK4nCgMKnLK4xas2xqjcLbM1s9stM+jfOUT0qNoKeO0z2c46WY1k5fNkL3Fd5ZZ1Zx6b96wl
m/02r4JlBTZ4NesQZDSEtNbwZdiI1ARhV25LUW2mGPTD1tMsFzc0ijob9vE8x1mAYWi7/qnZNWnS
CXJBchcW3KNAL84XW73PU7Ls7lFw4+c/5/NfSK7/+VZ3lb5O4Nio4gqdrD6zPG14vSbfhofbbwo4
EoXBlGFGKd4HFu6GuIUP0qyIz2EmMF8Xe7cubu5givy3H2K1kGklQoujcUE7m8KRP/HRroNPet9S
t4VNsLiZNmulwIjZPB3yYUIIKPrmrmiDvbs3ra6EtDJq7yGC75K+G/RjbC5FwIqapwiyc7J483AR
JQc9zQaCYc/TBUia8pzKhUG2wzaaVXUJawUkEOoze1+z3KfSriatUSVBYV3QnT9q5YIhgs7MlK0o
e/u+c6Fee/HG/OynRmRSLIdB3NtWfVNlAc8KWLH2g7rFfpTrTkJ49dzXdAHEhCqCjzh+z/mAJCtW
rgz0oUgFoz2lMbAKKxfnkPxheosSF2d/NZtwwMOXdcbb3URnl6u/Q2VFrSfNzSLg4azIOscO8C0M
En8sAqQ+iwbDp/JnW3IytIJaPN83/q16Bpn0xD4IVFRCoRXyu7sTUMKN4GvFZak6VwgK4Amv/BvG
g0o1SVdnFiV/S3xu01xQKJM3f8dhccYb1w73krN95s2pur0MACri/Sbz+93bkqchXCkGTrz1Ylpx
XddD86WfQVH6Fqi2xOb7VdzpKocM+TXhwKTVfSEinEBwK6PxF99YOUrVGeWgICsnODchWERkcr0u
x6AQL2nCQAUXgOoDIBNmupxZTeqTd7RBbFQPWTeRd3ZmSjJ7mpOs0l6mEF05DbP4HsMuLECJS1cd
UsBh7U9Skv9PyrMjg1IjakXnM0nYq+NGoWMVO2YgWPTAD+Ok2JCUjxSBrF6VxKXh6kmuTNMCkoBf
EJmHD3jiFxgq8SaPfjFW4BaDWoQQXKMzYVRfbC+FklL2523Fez4IPnIkoBvLhKzlQh0xLw5yiyVP
zU/aHKFctMrOYoOuSl+cOnO/b7Zea6l8QqB6uYb58dGGAMF0Ne3uOuwlQ6Og9b6sYZCQR6INLssO
sCUuNZxjhMCQFuncTEUc34tcW39H5ZPLDlE2guOuAaMoYRXWGcPTftP0yxNnmDnMGNimJuwPz2Td
qVTQBafGt8DK7iPYjOhajAAPBzhYfp9hxQgnSE7/fwwmcir8TaKfQk8fi+T6I+csoZrr2hwjuD8V
eozrFRWQ4IjzL+jJjlfvSbXmjbQa0OrSy/ZiA8+BaiBrJV0oFoywa+53xKbHNtRahq8HP5xTzY5q
q/MAgyBPbAUeP+6B0+2Wmf7//ZeiPw8FYfUb8U/CzTZf2AzVuEbVXCN2yOngGk8EX6S1Abta3CDF
gvj2dbjlXbTHUkFVNMGAu+oELM0I4Y7okGLENlkX22KgDV6Mk7/XSDzGpjeMlT/FP8yUqEUP/yls
rOot/vrewdm5DnxSfIwLxw/kGBMSQs8PqNNJhhjmJRUzJpiGYN1RiznUa5kG6xfUK1hgKHJZTsx7
ZxrYjQoIAWtR/0reWZ6neaqXxK3ixh1LIL/BeZfVuYMpr4vXFNrCBBfcu9FNtmDk6XgVTYa3rhf8
K6voQ9WaFr+2NazEab7vL7P59UtzlZ2rU+p6lWgDWgHoHN9jM3Wep1o/6n6fajeZD2++Fy2WIaeS
SrOIamA/MWLDEfpVcVBq2KK89b1bujFujPtFnNN/jCf8nOq/q+FCGWx96PcyNapmUTtW7ii+H2RJ
38H7mVOtmG4RIG3dbZKB8wwegjM8ZS9AYabWSp1LW9jxCtpijCrrYYD42l26ykNAux7eBPqzL8FO
iUd+7iE3GbV+H5itEkix3d3S0ZPGyFCychIA43MSw6KcNtBszbA5S+TGqxxFMQN5E9MtuV0WVy3J
AHDkimgLx1rO/wkCRHmAx+nJe6NP+fgU9Pp9HIWQsK32CU3h/+nfYgZofXfDaWHAFI2VR8mdVbN9
VCDYQIzVuBPrQB9RQUI1f/0ACU+jRKhkXBZNTIwV8ohA39eo6CYl2qeNLpIqppDeGOlxIErcUUKl
jylRrV9cKbrzFqTNG02Jha8ZUV9uHeBVv9PH8WHivt+BABwVpMaxt68SRKfpSoEvQaemIYl4DgTz
YkIva/8yraLnWKCVy/Aswrhfu5RQg4Jy4RDbEBiL6ULynN4D9foasRqrxw7hETXU3Szf2x4aUQEc
/Wnt/J9UJ0sivZ04IIb5QYtov/ZSWV1Kyj0lD+i14OtvuP586kzQGDXyfZN0T2d5hH22e+Xx6OA/
3vOeFQ8F1oIam0RCzgpWHy3g3MPnkHtaZuFxzIFVjrrR9AtBdxqKz+29oWxJ9w5tMkALnZmCd7QC
kskJkV5VLOI3pH0x9d08V/uCZwN8Z3Do1fW0X34J7uNKj0hKUwWS5Nl/BBD5SLbqEr2pfCj/uxmG
mTG6NeSk7fbVmdNBleIyPnD/cuU4+Vscc98WmoXeZyICOBIRNAWYYSgbiPGdzSCGQCLIorCrY7/m
9Wb8hB6gpeeeHE9tBudEeKIp1a5tZFWhJuGmtwteDKbDdd0oYx8QMUhuTeWwNdMwGrxFO3B8onup
Zs6kQaCMTe6JyCIotw69D8WNmWFpo7Cc8thBBgOU62+8EorYt9EyUXiWjqEGZgXQO5cJGOEiinRA
6/T+K+gg76QoiqgrrUP+Sb6008oCT6DHBMp0s8QH5XWbvw2qCjXWh6KRp34YkcCYDKyD8etKYE9G
uIRp8qXKn+M8lGbtC5byjbTa5k2a0vBbWKMC/h5ryuFuqEYOltQ9AITFJOUtNTR4eNih9LHRPwhP
EjzPK+FJuV5ElWsp2/7x44CczKZgxd2ds0Q4TYByzIJevZCjid7n+VcQefvbqMo+WX1WoyQX591h
zsBwPFe5UcEXJfOB/Y6gc51CGKBJQffSTMGGCunxj4aJmrpfPBPDodU0A3PEJX1FSfwDmvtHYe4K
0oIT4XilGcg3dqPwur0Zr5PVVDtMOl2UGGJWkc1sahm1wf4Lxs15eI8LBSlw1intA4d8b2f4R/mb
c7qnBdaknZiO3X2F4UnNxm0CpVME0amxLCfjFC06pThbtecVj+MVtF9IxREuUl03yhURFXygrezc
Je6C9FtMANCpwIuZHhv6jH/Ny/3gJ7EuLB2AhDW1b/sfFHH4teF0A/3SeaqE7u0B3y1RqCaVj1Y2
5PTpHWMA21UH9HD9RYgJQ5gcOKm8aw6J4znDQn8WTeW0xmiq1fNJgNw1sle8ewyzyBCh9AfGfED6
vfps6mLPli1xeEikCeobuXJnU0MH68ecWbMnGCucNuPaBLeskDjlR2EsiSsAVfW6GSlcCtI1l/3R
UuUAgAfU3CKNkDeGc36B2J3XwbWrHSj4gALrU/lplw5Hgzn6Olq6IF+IJz9PkmudPtcvLANQrdMr
LfCP5xanZYOTSJGoMvhdSdFlCH/TUvUv4gjN6nmNPfbgjcJqieV4w2HGbrHLgHRibWGmaReDTgBQ
Q2JTyMRtV/B3gl/j8YZ/uDGw72N1Tie3d4JWR/vV70uURSXJP4e/LGo01mEhZJAxDqaj6QDCxhMO
KI6BDl+9GNLz/ZvCvAVFkn9WF28sBa9hgesHAZZlu6kixJkAPNTrTIn81GFBd+soLdnk/INO+etI
QO9yI1XOE0Azrc3XchZp5BRTObOKFvv+E0UKLfMtC2WqJdwD8vQtSmlG7LKakg0HHma3UplXqcXH
ae0vpp1NpTp3sKPmhWw+GfsukQLi1KzdurMscDf7ClB09Ba5J7jSjpDM7tTEJE0ROisJxK7IfsNL
h+QNlD8iAg8aXBQ2T+Mv2xndbx+xv4N/2g07YTji/r803HFyqfjrDNTeQMKC+SHVjaO/+aAOLr4M
ST5D7ddgXgMwd+seyweJn6MSR6ksNy2Ggcpl1bt01i5Xk8o9jAiW7B2VYJ7YI0VKMJ8TiF1G5cUK
fz4fpGbrxCSxZhJjWne2VoxrzalB5lOO0iq5h4kpYczeE9LDlSnYlskOYcTdGOoHP76ET/RZ11r2
uCv0ZyEx2AS0FV7U+MZEz4L8LfQEkdpLj2yE8gnY+oKqsLh6hNYAq/c4YHuxYBloYEQcfcCWiqe/
UUV7+/GlH9xBve3xiDPVeFknfFSmq3n6CwhipfugiINds6uI8pCvp9c5hN9JZBaJCmFpVoKs9ocB
aNXSz1ADHQatqjsXLuQ06f9jXy5RCZJ3GhbSMwq4oBqRdZZWHaLdb7aebjcwL/0wNmI2d1ptMpLe
TsR2NRiuHfK2659q7XeQRrcr8hoWIwhfAvl+TXygYfIc5tvzJVu/inReC0paB9DE8GpKyELS4/23
QtpkbGmOo8cweI4e6Xg7ZDmSX9JXMXD7GBrFv5Z3yyOOL3umk6uDj6d0AeymBY4ShJZxT79Rqxzv
TeduxiBZBVDSsvB6kZbdyU4p/yzfMYEzwqGixEnTTpMZwWmkhyVWgf7LaoM4N3V1m9QNnKoK/mqb
I9zVhKcL8GjNP5rcxAKZaKaQ1ZPoDZLnuKWSFLFdZC1eicD9aL7QGe6cIlcHVGUhzGPQrtbeu+bg
jJfIx7PUGuJT9boRrhnC0lp1PXpv5b5YTF/2OLdebSesvbBD3JmKtBX2ERO2MOvv3Rww/kQ1Utfg
7ZyF9q39fGEtRHG2phFd/PYZbbL8DRfbvYuLvyy3h9O1z7ZoyX8xhyY/k2il/4oQzzhQAuVcwnJA
k33988jWmZH99q0VphLywE8T37XJeC550AQTpNYx8MSDQFvV6JjShGfX8f5kIvmCccQCcb21tRP6
kdOFA/Dcp6dw/ZeQdcjLUZeBWF6lb99FJCJpSfJoZHGT0Ro+FOC40KGVjluILNZ4V36wmMIXj0pA
kecjXyzuwF9hLwa7hx38VMPqvQENRdFtXu16ESqUVKR8TgjaZdu4hvNQz7aeCU2p3cxWUYeotFRR
YvU4+hmMFkNesjoLWEjNAdflEfpyIAcEncw9O2KkFGnQ7ArCQQ8NfiIxH+bn8KkarITw2drdRHvZ
kLjNW73w60SjzznQdsMjDwfLTC3QQXD7+eRiNTIKV5GHKXqewSFE8Ii1jDDhq5vZ/5lm7ziAC+fL
ox8HEhSFKAaWSi9sThQs4GpwKHrw1a/uNM7vD+hyqSWZ3A+K+AbI99A2MXneQ/JCSPCK3PJ68/cR
MKiW7ECpB/PPm8skJHrfL9Dlt7yMP62lDlcREl+QNQLqR3bD6jW17X3n78LaZcHtW7te+jzrPDUq
0DeSGqtEbFaI6QryN8V1IDfkV7MCEVgSYUA6oshNfFZscc1iToP4uAXrzzjf5tHAR+eIfabbVH2N
kGGUq5FFdm8Cf8OhR+UgIA63/1CGxjOR2rcsmaiFhuqbxnilWIPJskItZDcqQYW3/iWmZj2nz+Qc
QD4ItvZPoNlajYRnq1nRfBB/jl72l25LAUjewDBmGyAM19TSD+cV6DwX7EJmr2Mg5YGDTwS2D6ow
yUo59dxK/UOzJpxs9FV6DtLQ3pJGvnnKlx1gi5mWqt4VbUv3JFKJqRALkWtAC0r1Od76sMppI09o
iHwlwqmM9LYawUVtIbi13Ho3RsfgduTBMLOQBC2x0Az2kR8p2EfC7mvFIrFcCtrdpLtp5vnD8N5t
tP9RXkCIgvNcNJhx3wDgumguxYmydTe3SeL4KlafkDCpRs0vwUeUww5SVnXvZH8KgPbNrS5bkByR
0BDW1AjE1qLCqVvJ2IdSIgEqEIQLj6W7PHBUYrcJKWbTrwBMWoRQX/FD6MMkR/Y3cjR6r/f1v/KM
4/SfbywTW92n1Ioewb8H4bmY+depD/UBrew9TEX+BSgKSpBahtEHLEXITSjbqmasJyRlIkG4rp8l
zsuHVuYa6RipnECw37x8mOl+chhEH2blu9ipftv5BFm1rLpWYBMxBAjuD3qxhnaiCfmR2YPDzph5
UuUCohOfSu867jdXRbzN/Eh1GICCVgvzi2UtZCXPjFH2SUVVFRiBTa5hiC9zgVMICC13CS0T3hTo
KUbc2JlZLr199WWBxzEwWT6jL/KHBGO7EmAIjxap1E7LHTLiLCBCT3ugd/VnM6E8/hDZvyaPRlFD
dqBYHh/Kou/E/yj8B+nNfLjMRvFm2BMQJywEJSHfZd70Q3TpZSdQefc1UOpr2TmK1kDamiiBi7uh
Fsm1sPmMLchFnGSZsNTe5IObaidr7EIgwopx43ScDmnRjZtdfi9yYS9/H9RT7ZPMwt6doM7g5hN/
kLno3J94Bdb3j8zV3ibdHmRm62W6hmwLRZkYZCq3DpvCUu4cfjXFuaUVWAYaHbd5FlnMumgy2TYw
N/8AoqkFNbeCNZP9hYe0bckahPnrX3IkZx5BvGuxcrNgmYLgyeCksZoIAGqIywidBprfIPnloqo5
SpEdVJxJGFQad/cCVuiDqfSN1rNdYPly1TkDZqCxdNL0GDaHYl9wTR/6HFn/EHC0niGqjsmQVOb5
7pZnGOTRiOr7AKjJWT4C4NN6z7XK/VnNAsN6mODR28vJ9s4cjGAVU6y/ljlsAefw9/ccFh44mYvH
QvZw9QTEnM4Urmaahy0pNOSsFbzzXCGmguNgao2Rv0PVrUkXV2VAakrkE8tXDVHiiJTU2zsxB76Y
irzUL70H9PBKXidLqqjbviGiusgBILZywHqfl9Edr0uegCOc1bWbbOJo2HjsqaTLUsI7rH6L6+8q
EZ8aFdwmoEjGJ486maRwF3E59sHX7DkRFZP1uIHv6qonFePIR6fJG3arEJtc3xmR07TFmFhdoJt6
z5Iw1iY9xuGXcg9Z7Xfa93PDoDtQAznr1dmJbSvsBJj2EwT4bqZbmtOHTul5Efcxq/j++Lp51DxU
DPNv83/AP3+zWC/DAGBMVTxM67yu3tavKQaJ1jKDnrVdL1MN9aGt8sKqbtlOqB7kIijlPfGmQ3We
h7uQkjsRi665BR0euMGG+QFdQw0JLexxRHM3XLahm/HPwNEd/IPNxkp1nUvsAcrAaN+o5Rn9LCqM
fbnmwtcbyGGYIdsVeU46pidIpUWpIJaCoy0fpko6v0zfcdprQxK8GJr/gHyfHzKnXdBxmVx4Pjxt
2SQ92lgCUB1CuQSs0KSZoMcbnLi/6SroNYwMlz4KxkIvpBAU/d8hf+kyQjrI+s/1mVduZEQDUdNV
9Xc4J5+ShzEATzpBukAUPHvAlXwo1gH3rUvySSkk04nd8MU4h6M9spq858yaVEfnfU3Ct7Ty9e6H
z8wKflY9yOe7PfMhXmHqitzryFKGHr1vkvkvgxoulf5gwFnCgDyqy7p1wDig/aU6Zt0HodNfvTGG
nJV7fjap5xKaQP2tU3SJrAdlfgAuExK2knx+FD81gqKoowcbxBkp5HvmfIfeW6eD3xmne9UceiKv
jDWXCjwDoMy2iAo60A5dXWRNjsg8eqPfD3XT33/YCEBKds3Uor3HQQ6bvhhSvy11INilWqkcLqWQ
tG5bZDnP1CWvB3FbYvsuTmLQ80fmCTRENnr0VVc7VSW/SuTpaB179xVheJVwcgD0bKzxjijhhakX
zCoj2gWc0NMwXInH7Y4cU9fY7XamoC5qGc7oBcv66Xt/7xhE433TTuif4xTBS4+hswyK7LlYD8Kc
4EwAqGVWiyLVNnKiZ7NDoPBOHTT17o8z2iunqevSNF4J0dmTEoGKzXNRcvtZ984MAsRR6PKg3q7t
CbxcaQ5ht8F8B4sIcZSDpQeHXGrS5h4dyoUArqfi61cz+pmriJBRG+VTJS00s6UJeBPXvsJDIih6
KMfoN29Wfdv7rFJLCm4RRxUzqpeEckJd0Odcthj/Lx2IskfKQb8ab3Vdq1a4egHiPfs3cIjYToO5
g+uXMC/DdXHEipIz9NXXILaJfCCJhQqHCpi6fWhugZWce7LgfC9beCYOJ1thEQHSisgUrRokyyyk
NQkMegoFvfEimtdgi+TU9nWsSlTrkp6Nl+uUcdQaT+CpjXUUfHRkMt5ta6h58M/LbOPKIaRqftzd
MXSTe6PZk113oY2Fau9Ih5xvWzfuQC8vJJhBdp820PS8pOw1riWBTqcsmDWDfw+hq2zT7RkLt8Na
q9GTzgJxZBoiSzEjOKhXBzplzZ/yXRvb0o7h59VD5ONF8UWWDaGjQgS7mfHn1Vyv13yfYqW3mlf5
sBlHry95r8VQZVzyCa8IzyRb7/Bl1GRopUbbYaM1QmUc6mVjoKqIR4bRZEEcrYFGGbvlv85++2QX
FQlNjg+0YauVVwkWl9TVcHKejM1Hm2SvslaE7Y6lZ/fsBFp6iPScBSELcevZA7nASxHrY5fUBWPE
2F3/k4/L5EMjSjPWbaZZ7bWu5+iz6dkO5WQgIbhdKNRR3NNIya/Ss3KlOM6UYLrRY7XLSQdYyHgr
fu20NOQdBpeyBfjJI/Sv237MsVKARTLLiMOUq1KGOMB7pwJkCy3+V/1etQ9Mjfo9jpY0R8npk9Ms
bmuyxHPzjrjLtB9IjTDjC3a2EtZE1y1F3yF/o3uAJzr7G+lN9wRfBQ3VoG6sZKt6JVurLorDZQ+t
2TfDM2v/WBaMv7/zO8hNv0FgMhRCYslvcIUoXxot2C3i+nzUdGwnSfJTcFOca5GTL8kWL6q8TqnQ
OzE+gNe1RH/kt3yEHBDth9j9TunOz9M4Ec3yOdUwHLffcsT4btUvHaIZTpQ/iTTYrUW9A9FMR7wC
F/WK1KTq8gozkPuNVziBWkGA7s482nUdxxdFQmToyNwPdF60h9eefc22Lbl72gePhsdAnV6GgX4T
VP8/bdN4xbmd8xPEySSNlGVzroxu5abdw/UK+ikvRFvVW7Gd4/ua5n191rMp+UJOpc1+30N5s93V
HrzGSqywRYRgmWCyag6Etxb3J6URvenn8Uybeiy5Fc2E7AhS4yM6x4ZWjCca4ywx+LjVgz9YHyPr
q2SmrqS9OUw/8NUmQZW3+0hBPpQEBohXXEHDqY1tZtVhaZIDhB9Nkw+oGfgnzdYEZ7kr0HH3Jr1d
DDY4CgvQos+FrOvWf5MOAsCZU+yAo4b5YGsyP6RBXBe9lVHtSrG6PEuYN8kMyR6NuqMfETWfvjl8
8iEeWpsHtRiilpqv7N6pWApglzLGODE+h2eMo6fulWMx0SUP9a2cvo1SiYj9EXLqYjUaHV67Wu21
9+v7kzYVJ/6GCY68NVAh7WW+g2L/DPwVPsG/UrTAtfCz7W6lGd5jUjzGDV1JOc+AK6T6zw9nzzsJ
dol75GrFtDjCqyYO6E+r1y8mxNGINEvE7TDjucQTGL20aqOC1RJnkYMGIA1ouLyccU1+qNDtqcx5
TxsY7mBYCt6UhCyRUd2wFY6vfxgx8GsyODzgFdrDUaGSpD5RJS45T3Bjd6kEcEYAATqDLC73zGsi
bQK6BN7mYQcJlOpqxJcJElfaLB7hJggd88eSvOLbegDUG0oKSWRS+MbWva+HlPccWrc7Rwg8Gfef
6jg17EuB7DFMyyOKLnHJ4yB3mi+padFpLj/EA/5lLhSMTrzu8SggDGIfRkPV4jjxigKH6+ZNUQv2
IKbUl0FtE52+tOg/GKaUg4oGsRo5qH3/J6zx3kssTOPWYkwEgTkt0LCRvIk9Dv4frjyEui/1VaDZ
drikkUq/Cc+wK40QuMMIesHgTz4qxAkATxCfP5oq+vEgFrhnUfxMgcovWZBCJotVzY4kmG0kyEUN
2Kaggkr3JeCiYxE7eskpFDIXxUSh6vZwf4M/PCbw/lLIYeUA6qLC4/N/ueuadQyokltbE7TUX8zq
CFruD9959hPnBBnTIvIv/TXOgI9i5JOxzGSdTgxvbSJbDDMmtr2eMgoYpL2kdkxopSr8kLW4XSC0
huT6XCMc+v6vuoj+s+g8OrNYm1dbYoQXcDSjm2/FtTjmhMlO+qlMgwgFV1js1dg0w428qgImYJO3
toRc9ySXG0oOraQO4EnQpFCgHkQF2FGlHE5wWJYuEm4NU9Zr5x9tZ0xO2sNR2h6DiEfKBIOXgVy7
Nh1WQ5RvBjcXHeXlvww/LQeaSNeheWrq1y6TtQbLWNmMLkc1drBB1q+OHnmocSzcH6wWtsIOJP23
5W3fejX95kAnTFW+Da2Uu6zAXSXr7XbVrpZcBXco5xb8wOXlxLK7olQFu04vAj60HNZs0BlM05KD
kSI19EuzgV3T3fdjEv97fe0Uu4WJHmRlPJ01sNPO7lWA0hAcMR0OjbV7qEbu0usEMT931isNVw2+
TGAEfpC8ptk3TB8mTgqRSZLC8o13v19Ix+BVJ16Hwf53ZyOeLlpUiLYEP4mcy1SJr4pB9rPxE0C1
Nn3Ss1d3rIjyfwmlrZn86qFe2OcZxYbbYlqRyzSoqPNEHqDgqs0QAWYntnkETkSis4kHQnsu/KJ0
sl3IHFpp3aU2rQJoUfsbBys9WB5vVK2yXadGfSw69F//j00tU88WFQkCbEM+hRHCrj9t7BBqPKf/
nWotG3bnGCir7AY/dQ6F8/UI0exUmIsf9/RN7oH7UmQAETHVqLI4DVNc9KyVHt2AN1oBihKlX4AJ
n7rs4AzEVuomdyB0peuZ6f6pGGerUhLNaABzDwnsGQlo0gseNKcUMqgeFSf+PFfGjETG51pGlRcW
doVhhQfU67sobohL7eAsUsfHV156qnqBAE3YFExoH9eOgMmN+RIp9MlwKFKlUlvTERVRHokXZrOQ
3Lp+YgmdZqCRMiGbJmfyPY3iZZwPTm1fwtjr/3bT4TGLWoTN+tL+KERcuje1qWxZ+syOq/cFTwGk
PqI/12EcyK59Ls/kLn1gb/PwCoV0ZJlUFVfgK7NqznpKqLKJnnNWRTb80FkvwBEdXnIwGYbYMawt
3iJ5kpZJexeHogkf4ki7LLs+hUdQwESK9+URPd+o06BPKLDj47VrqEgBwqD25HhWF6ZWI7+beqj2
bsBvKqSWiog+C8CIB+hXW8nnmUPQhD5CyXD8LPZ1fJeoDwozJkhwZpEEKMNv0KLXYmuQAzAF1cft
o0m7utpxpZYOKsnAFOrlHG0pD/Y7vWDfj+3LfGvlxDzCLoY+rixaUL93dhiGrt3Ikp5pjrmofu29
Mf/yinS4ZturacuZyXabnFZCrNrOGw+w0YvsqPBvlzcBe9hUOm79JNgkg+PTCjpifJMxbJkmpkW9
498sdvnIjvdGuCuHqMmRFXw5+whftQm6QKDNO/L8cUgpp7F3zZk3jc7A6y7dTWCX5TZOageqwEAT
qpNBMCf3lzkOfCy3N8FU2kUslhp4pyayJXUv5B9C5WsrQUc2738WOjsL/cLGO9ZAM89oWfUi56G8
Q0obwswmMpU9/2Bujq6tRBVPoIXOBp6yLuggH+a60FY0SGhWWxTe0EPxPV9b0jPWnQ06spyrDNNI
dEfuepwDRLcmTQ7pRnuarmdLtHoypvYxn4yBgmDqiEJsdvZ11w87/hH7UFb0NtXIs249T7TTayKO
Ctw2XmUO1ZG4GGC8UQ/8eD7o8xaTOg9LpNBZh5qGJZs/laeTySzpXyC+tfOGrjz8+ruylqOSGUl0
xBYqn45HBcK2vmudSeKv3spwqKUKMHOCARjbQ8q6wBlxlyN5cVPmeb/uQaUONdG3fyzWMUHeepiM
wgVXWD7mlwUUygVJilc9F2n1rXYdYsBm75xjG1WMldmr23NcFUXwFFk7YNjqQkR2+9kuMvmOygpr
U0SBt2InTjjnaEgo6Yb4YbBxknCo+ALG/V0VPTzYs/VU3Hpyu4JjJPgNjmDMsBFM8RO90X0/JTbX
2eA2UeqDuIqrm9kuUt3h7s8ngAf3AIEn0p2Xoda3b0Ukj63EDEMJOKdKNIghXJWIlxDj0nZ3GHFp
+hvWcRbEkUBenmONmqDLuM6ebKUQXOWeu+MqSZ6TrH+Thp8RRVYJwhpgA8DcpAvwQoFZ7EkTQwS+
LIL3QYzjoLSy28rqACPmMKFeSkm+olZLIC0GYi8QvUHIEJf9SEFvllg6IPwDLeT67iN5FeOtNqqU
ghgo7tJewuPxO9OHRICv6Ja+jV55hlp9WL8qCuL/tIDIfnQhFzK0jvyf9rITTPhUtA0b1MbbyWMa
Vh+75BKJ6C6aI/kEIXz/16AJdg/VNEAWN4Jd4T5cm8PGIbfz13H4Erqy9VJr74v50CI37a5FKR/7
DwQwDGZKqdMg4oIBjeIRV0LhFfaa23r83rsrYPg76IOp9vfiK2/8fbaliJJ5n3c5TJJYN52gOlD1
Roes4aH+B4bnKctQCsfqbbBin4CsU4VtSLIPEthqkfnHRKneQ2JaBCrDs3CNxQ9r1QblITYCR6zF
Rq1EHb7iVsspHAIVMLhTO++zakjGNMthW4vekgzTk4L8NX7eNSkr+BkTg7lu03uLwuXCsx46LivL
AmuxzN2p0K3NenzKqQbsoMMplkBVVtrGMElmwnR5YIBLKcQZL7xv/knNW5pvj54/FnBXOTraq0JT
juJDrvyH+1m0C/sjHHhyT0sxDjVHcXlFU6cBYcEwUYi353SiE6cEQzIt+ZqH4TNLuYvOHm21r8/a
+seClm2YFFa1pPiQzJXwntKACsCPNW5hirUounxEujEsDNuP+e29trvNvkHf8hjhp+BjpIcYUQwa
jbseIZWfXv4aG3HLhtRQdyezzpsC0BZj9hut2XxoBBmozGMQMhJSujgp0LpSwBfqvF5yg9y/Ouwg
I3/PlcdkSUlIl7XGf2mAu6/M0QdUiCIRNjl8Z6xT5iRQt2xYbqfMxBkaipjRIg/3v6t/qnecK1tA
FNN9DfS60nA2biwKutEcKmgQ/4AFR19Tk5tQWmV0zMnnhtP51dRP/xPS8Os0abdbOwtiJWh5bEto
zYSSwf9M9NgN6BfY1MJiFVm2LpgvMjROxkw93DZH3ujmeIOLXVgPSG5PEtLQv3wM77DXddAEiy5k
S40lGbr5ZuDNzR0s1Cmz3yL8lazEI6JURRijn+yHh+Zv/FTNiEmMBOWYx1KgYOcIvqqvkC1HV9Gy
YScHOw7ODb8/Y8pN825V2mvSizY2yOxoKlSKrAYyR+mUBG9LYPCMkKajiup3HWhobimvO+/gtCfC
poThjeT5BLv5Wc0MWw4RYQ6ePOiLLGgkIEQWDmT5JD6WF0AXbprgXXtA4EcZB+7R/9Vk7M8L9973
H/YIu/dtG/PN/i5gKY8S7JW8//7PuIdMrRocpoJ+EqZJepec/07CjupL0e99SOcFxoqhshSM+pQP
pG/TI+Qfbm+EOCAXHhAzd4t9d131osfCnWBZZ3Qs0bECEd10bW5tWJR+T/2NQEM/Rm6mCPHfyugt
ALU4LEK425cJ97awvo6hXQEva4bp6DgRSGkUdCqYk6sQE0eLnCVsVC6ZvH1vbuqYsWPg4YrUY0Cp
WkC5z9OfGK+gP113KntUetEdM7eEjJnPFWB8XC2kmoQeUMvLZ/c30aQCxw8slc4FIq2XVG5MfsMV
OYWP5aK23vV6/2O7QTe2yloRE93OjWGjQHpPdiTa1cVmXnjPsi08qY4tIv35a3H1fsvWDvDl2Zo5
aRIOQx0QzwFP5bEtptn7wNahRjupsvQHZyi5VyyKS5LlrfSHHUvz6PCQKwxMkASklS1P8PRUvrLd
pxMbTBhmGHShW+2TVvFH5WkF8kgYBNjDcWkFp3lX67x2Qu3DaHzWJxgNihGniafMbSw6TL4yf3x0
Cn4vrUOeCbiiDAE6FySEYxLUWlXV6bcGSUqp6XrxxKOeRLDFg1zrDVLM0uy+eblUkWXKqZ3dbJ4R
N2ddGl5eMxtVbn4kcX3+nC+VLaCqaTNlf6TrWcNPW3TPOS7GI/xoyylvv67rfux36QxQyIdIuVm6
VlzVmldKultu/syMjmqHwN5G21298rsU9XonQuQNG8/1lxocWHUShR/5DfTH5yNlfL8ufx4LfTvA
Ll+pYKi5DdWVI/1hn5QLToAPLhpp4z8SXlrsPtI6cnXtTWiqSZ3Kl151cX5PdHD962BHc0RrwFjL
y9qSWL4wJJjAyalc1TLFFDr2FiIDp4cA8Jlvl8Yy8Wd30JjT2UjnFUVCnRBV5C374Lrac4E95Qcd
3QcnHcqSJLGwmPApZfWd3iy70SRzWt+gQHBc/dVw7V+T/kzYbsbEvlB9xubZcrU86Bru23BAKgRV
PNWyaUpITPUn1MqWV21tV7hY9mLlNPOrqrjKArlYxJ/VYbT7v3A4W83JMT++ppILYksyxryaOmuy
cImBVDoy5Nv2dQesH3Mv9fMOGJmnJ1mHhkR5mOalBBtCTVaON0LEBXUytiV9EplPpDI8+UsvhhhA
iAzbdMLbNxOaIPJDv0ub+QnShtT70YpBCDXbRgLS/vOswS4RwGpzhGn+qvEyEF1Uu2KPB4dZu/SL
tCV85IyS8LZ925IlmvncXEu3WiLHMa8qTvtlMlVqM15kVYasfVwfDjUEqifCblK90Y4W+R10mlzc
3RdfHfJYehYZ6GSOkTeGq86SeFoc3RglStvXHq4W3okAAUyuKGFrAnh48LiewwKPngwWq7MeSROH
24qbc4i8p5FaujnzSD4ckzu662E7pDL6o/XF+ccaK1YdE5PfJq8/8Bru+FEKc0NJBuI1djqs7Vff
X8Wv7VToei+LC/paJbypCRGlVaLzcDIPE8vx7K+pQcKb7ReQqDFcjmHyUSSF8P9CWCyyNJwCq6lo
3vG6KHPKnA9/CirEGJixqMfu/2uM7ovCdQoRgT0xG1YSbqP/7aG8aGzy1A7E6yQivw3+Kl+PZ6fl
75LLuE2akxr3c/GJfZYfGODWYX19CUFqm8NtwXuONyoPM8Yldq3e2cZN2vPG9+NMXpFdnpXKx58k
mWCTJV61ttdKHbMLJnek+quRLG698QxXjgYjq1F6YgJngNPzaP3pac/9g2x22f5ZSBRjL6JS6sux
3UMXzm5vGo5HrXXJKZf7eHSC5UIu0brxzUaHLWhxznuvtpVraKN/iGrkY7NwWFoU7S2Uimz33pWh
oxjJsFHMco+0bAYDrZcdiBckO9qPHS+Xq/8klgaFfFWoq5TQ/gxnZwNCwZKAsPHBtA9j52eBkQjP
c7+StNaZTMqELrQhg3qLETh7QkV2lfXmmVy7dYjYCzLIWrTSXLteJ1aOGpbU59uiYx8FxImuslQe
qtsukdUl1chYPPoSEu+osWvXbSrPe0h6Oawct3sPZXFB0pUHSxTQc3ty+VMbNLZdk1C0Hj4bLoL9
Kl1QSdAgqMSXv4N0rn3FmUFf3WNX7nuRFmMY8U7KF3w+Lxcudrv8JPV8uYIjFO55iSjj2PSfKUJP
MYny01Hyne402DPbOXj3L2LbFs3na0OqX2G9ebDYLN/8X27Hh5ZWznx4BfuM0XofgXLb71mznO3X
ooFqsgjSGDS8QaBg7kB2f7AMBvS7RL4FfOFFrIg+5l1AUEb4MEdDjL4bxS/wIORXVHeV9ZtJjgfr
ktYOvKZEQcohbSymfpBxqeSDqTQaJhl4tmSiL5DUsrqWO9n2DFamGCCkW6hZgpxCGoruiOiMgtU7
VGXkDchZSo26DAqUkll02FnimIZkzBg1ACC8gJDEdgtlgdYSrX10aIPEq9+r9J1jioyAxg3AWa80
xZxuEnEH6pVFIseU5GZyU9c9JOswVq8aUVRvJzS2IFQi4zimF7eh1jLJFg3sm9RISsmcatTJhZKa
E0pB68kxydjvr+1gAtb7M/4NwYCowyodbERTWCI7hWeCoTrq27AwW3YktnOWR81wD73dzCABGLGj
CPgDedfDt7+tZhS/DU5ncYXY88kH5ceTDwVbKsuyNi9eMBvAHPLOTilXWtwFH8HMv+4jYghgcD5U
CdMbEVWttdtMbWDlp7pGGIIhJal+0QcrsutjGjv91ALI4GUWynQV46zavIh4CbKejCJgLx6VCSoK
wiWx0g3EW5szF8cgpy8UJIY5BJg9elwTDvf3uI6BWZTZlnPBQai1lp76fJQLD9heMpRujwyxYHN2
5VA08884Oc9sSUCtJdJC4GzZpwNuH6BolY351J1EsmHrS/UnNxG6r1u3LPUw2+JCFWYzorsnfrXT
LNHzMysnc1n2+HXTjGNDQ6V8j4JBOtzADM7k06/yl4SVzWsPe1LTrMzZyuw34t6f4Uvw+8CdZeFv
E6iniJGYwRYIpNibUpxBlqtUmiIA9A4KStsMbaNEmCvNIXALxlvH1OdFQWMK6mtfweNcPXiL80cE
bEfbaIZv9VmvRPXhBuOod2ee+mKKBeUjGFl5sGxwqn14YiLmNGM5jAON5vEztvGCmtSe8HXb7hnx
QIj9u9uC2tlqXF8dYGsanlS6ucjKz0DNh+c6fSBmCSwAj/DExuZcfVx1BmV1n7AKyBYd/Rgf18NZ
D5AbZmf4e5jeEUlmY0APS7n4qDcAlqguHqYyqQw8sUoSQO1Htqej210xwI+/gHFLGQtLAGnHb+wc
ctzIc7wDoZQuqGxSkq7wTu0pWhgs1rigzgSKm+49NsDF7FKIUOFm7qOBKk8hnCjoA5Mmon/kFXbt
BmOAxNrngXp/Am1Rdfl9ue0B6BtvPEVnlycGv3oBwij/Q915g5+JVwBtuSjMG/j3+WntBGAfd6oL
NRBSZxSMGW7758FdKrcpqP8JpAtVdSd+QIxvJ/mJF1cZHRSrS/glOOaB7dgEhow+7EKddZeuf8Dd
OBE2bei3dnprS6DhNYJjKEhmy551Q9bCRmDClHp0ac14qEywRAPxJUf0eYqV8V6lOz/knwxQJCxi
4C8qt7quteXFAWECsoXRTelTL/7sszUuXVzllxeWQt8f7i+WWmyve+GOsrRMENvqshCnzV+cFGAN
n713nFuLwshUzI9YE9U0jTYhxOgnAPufyEmZC+A7f3ffZqxrsvSIjBE6QI+YgEae59AiXNi2YoOu
oUB25k+iJTs5D0JmqDUrEMBM9P4aM37rRWK43Hq7tUCeL8cDLMBQMZNl9Edt2PZmhRu3VxK8zj0k
JsbWaXui2q2tMnvGGyQgV6+759hG/bxfQ86GWDZ8tIxHNvK8npSIMYIfu/d9MQGi3t+FwYo7D7HO
3QvlnCZwgRgO0va24mGYqtxPsAPBGimet0T94Z+7nnECTea3AnIt0BaxDUooIBojPRUMxDhOy3Nv
CMKG0FfcgSa8Rxk2y85PCr9xMEFAYR86+KkIMJSuaM8ErGylX5of6oqvw0uMEBZIjhqKkfORJHPr
rEsvczE9RA3Zxf+/ErCJeTRCoau8WVQmXKR6WIUDZMRMxbbwDfR88MvCSOd4HVmiiXp9JtsdHEuS
NKur/px+lg8SKYl+aB98xEKvzGOzaOjsfEdMfNwUCz0i74jGCGla0z2WGg+2GkLnRcSF/14B9rW5
V8yk6ri6/EPdixc9d55hW7he9Vm9Qrf/KR19z/HR9FxmsXbQNJKYVdvC5SCQXiEyFK6IokenSPYC
AL1iQyuu8REubOi4sT8IQ47Grw4UlcMrI96PfyZhCQfp7l+Hlw8fcxNk+IMARGEkQ2mJTFtutOYD
C+u+5WtgD7xM2E/rpfJuoGNfcTpfzXhC6xRXoDjwrvJLY35/qHzP0DBVuRCnv8txjxvdgqRCCp6G
8aUjO8V0uhvzuBvgYT2NsAMAKAJXlIe+V/twj4i38GUnlOGeep4Ka0T4mLE2FmXlTnJMjxyEizKj
7E1brqVk2AdHTP5KZUiBugHDgzNz2ARYPk1Noo5xocWEkCynMVZeSMG5oF4205UImIUx3a3HuEoj
YLeZbhdzpC7beLcU2CnVgaT+zyshQ2g+jKX5DObja4tECPgAuImN0QVzdeHrS+GOiUQ6XW58QR37
isPpAhttmN/439pUhg5dlgyPZe8e0cNBnBlPpxa89NQsndENBow4VJ0LeKgnbCy7OQHAX8wsJP3B
DwKAbUh/ETJon5+4P2kuD7Q+Y1gVCyvn3cdNXxDpRJRuwOrD/UM68mKkCZh2djyqVP/9GpRifbQz
K82IjndC2dehJesz39BUytK7/VNr7Dv0MuKik/3E+yaESdyJhHXvKt3FY9qei2qZelrRBL6UyGUz
PFlmoo5IgnDmzb6f6huF2bxInxQXWwZwmetz/j2IGVWRrCkdjfWTOkmIN8Yj5oVA4Dd+9TsKWGdL
XnvvKAymY1SMHc2g8MzhCMUZRuCO6WFaeszXVo2VvYPEqcGMXhdVvzv2lTRwYpHiiR9qgM6oqQff
hx4sNA0A/stI6OrQ7sW1MRYvRliIWcFZ/mlHMPdSlLas8N5iA6hqvwgjcF/iiA1O7p0gmvm1eII9
7tLF3ai0Z0Ko+p3v/95faZJ7R+U+Jbf8VYAO3eafKyCxtcpPf2Sb20AtX9UoTRSZMGpO6A3GmIQ5
kG1FTr+OG3QJddm9pxzi8k5fEEJgMqOxq/VXk+6bktwDQ1jC21xid4UA1uaJ1kSI03m4cnqFW5C9
LDrUdUxw34VpFY/wHLqduQBz0w7KNmn/va+y4QcmazjqrtUHWZYfEE2psM6kRXPe+TFUtdaUtHR0
ppLPJcjHt/OiUEBrb77RUkL8WrzGu5eVMBMPxE006+mLl/7ynjS5GCqQpGU6kr+orP4z2JfVHSUT
6sG12rUbg8RvUacWCThXmfXno781guRl+X1CmUNYiSxYJyFwNw1aqR3tMV0choTjeJOBcMyfAc7W
YCpsmdRtE9VV5iuTAIUTkzOveLn0T24HM8GDZXazgBOZL0rE8yrHuyiRj/KHeo8Q2oNjhqj8Z5WC
C87C4xBW1aZJtbDNApTuznA/XnPCYAGgAdYmjCL13zvV6abUbWprmhBjjRYlCt6d41nwlVtapceS
0ZJmQBWcIeZw6aTSmpve3dp8kkD+Gx42HJJEiOG4ocbDHndIArKkGv0Bx3qtO3Mhz6lgKBHB9Y8q
1IMBL8qXuXy9Hkh2BmPOGqmYRgXWW8TrbhZlWfBjBOGjblIh6bQ/3KupWyTI830yjGuP9Vgng/o7
+YvjrpSl+sGmAaymy31SHlff6LGhnYiSYrOvOZY2OQza4/s8PZNDQuFi4oKw3IuTGyHkfdBZ//T/
54ERtT6OQ8oKHzAslzCrIitNr3HIyc9JuBsqhx5TctbFdnqW0wJ29ojVdL/r8JYCKzZSIyAOTNMT
YWtobZvQMg9X54CHHnwlPwIHRFX14fbJbKr7VOsEnAuhfYEYhJG+nsxLr2nFda1RMT5kP84hqX0m
DZbip7MWwohugkBv0tpb3R/uSbgHGDI4bmmCa7H4Nx4oBtLfdlpe+LBZpa1GmDsyve4OyiY6nXWH
3BKmUmJ40w6OWMBY5zr8OT8T3jg/7l9oaTIvc8OHDVY4hx3OWqcAr3h+PsxXbR3Q7dqXSZzHAHKA
HKyem5ZycekHRd8DMFFOydsNitmOm9uDNUr07sKtwka8YnqL1jPKPeJP4AtQfXGDuXctThcRJnZN
DjTyurtzgns4md2Z6p9bjeJYqLtGrD5Ig9yWxJ+tCqONqeV3n/hKxm+smsWnj18ibP1pAnOpvNx2
BykqIy8cpgMMyb2RXBVtj4quHpKGAgmOCYgSVCHQgxCSjOL9HPZMsJ8LnYnCr+dQXidDuV5/T4tM
YHuZClKFJSYxVn0etukCE7FdQdHCOzuw3P/92ttX+XN9I/p0GvTjz6YEeRoDSQHmxY81SCXezFMk
RBulVKq2eiPQyaCNm+O0BPGI5h76giAIQwRw3z9LR3/Iu1kivKCgQf8h7Xh48LlzB+t/MTE5/Hlr
aSR2uAtdiOw3Ub/4sbYjn6iWEvx1Yxybh7jSKsn18vJnRPInkllbdf2fgHRvOqkBtUDURS6LcocZ
wN0nIzHLC4VCyi4NhCNsPGNv+irmIJOQiS1XphOm5XdCMduYLwZl+XMtKjwKF/yBcGv5zQVo/KeN
kNiQkBSJMemIff3ok9TAEQYBwUg4bxcjpoJtCXQ3vSH5nw4gbo4GbvGq/dZrBCorpJld2XhZN7Ji
Tc3yNHMl2Zw4vGuYqoGto4DpD6E1fULRqhceHJ+T0PImsIEX2Dd+BMSrcZM5UYGpPFgLjdBfOYNJ
CsDUrAkcc0Pmh+GY04grENXVNTnNY9k5Whykxnsc72DCmmJ8sGpFZIXSIr7lTopl3h/YazKDwO+r
UmciE87F25s+o5tFLrp192vBhoi4KQchtRDs1DfyP7eknFaATk4vNpskH26bFbg4SJ6IgmSfFk4n
8X7yXwdr3j38G/jeXjFj6Asjk+52IDFqUppmcTlZt0MzpCUpmRdlq7E4pvADeGFpsDWag4YtJfJW
nfYGmRlfjhkIKNhX0d/0tMKae4K9NFGg25tcEG6WtBle0v/rFnF7c8SBf7l95+14Nu+EBGaO4jnd
6V4mjLgbHxkYHeHkbwEjulvMTZhtApB/k6XCKQ+QZvgWEMZR289IGJe8KtFzBTZgOxoTBoTA6MH/
oJv7K3LeFCXtCy7PcTJMyUtAT8rhnPWjC7TQvRcvXvrUlfAE9XXer8p80L7NGF4l7bfqvJjDVM1n
SUjLuvVztxjC4rH5owH4ET3vzvJv0AGihPpK6PABsMmWa4TlKVwmIcPKQshcsQQl7Ppk4sqppqlN
PrDay+JndysOrPwcQBOyLfiy4hOctRxg2q28BanuBPJ1No1oJAe7m/W43fCMEVDyOT3E1nnWunUn
r77LO0bRxjbpkof/CaNbOKzQCW8i61EXoqD+/eV8klLCWVRZdabZf/4Okcghc3+psw/3Ybb0NNi5
kRXQeAgp/ohDjT8bE0PNfp86gzXEhOvSlR/+sQoX9quWO7VyZwjDNTuDkXxW3/74gTcdngoramDJ
R3HjzhSK1TEXXpaQMeHJlaICbQajWAJfIE9Uxgu8vn55cBCVERfOg9xt5jp/PSmE9DXVoI3hT3nL
A34CgLRWnEraTeRr/NcduSEgKhEUdRx6gU/moG8lVra4u59qtlvA1X79++sp+ALkLTLpzDZpFDY9
RuLar6eHwu+OXp3CvUB2a6Rb5S5q3+W+tJaVkHYSb0c27EqrPqoXGNbaEEC4Bv7anWAfupU/ryqj
in9eVm0MnY2gT6aQ1Lr2+OpQJjCpU6k68W91TIp4mHJRns5sGkWRO5ihCbCkUOpCrQxVqvGnPlMO
2lMFe4wMrn+tpnQqVEdQ5a+TTHsJOMNc9/9c/qjZTp1spKAU430uEwuoe6D+HVfuc1oihKKiHfIX
8TRT/aFdmvEbjkfZbcjrNVEMp6cQ/n4KzPhZZYWK77FbP3HUFNms6Lkq7slGbhPyKrajbWH2SzIw
pfpSGE90OapC3snD1NAWxqzhjNat1s1j5kBRL4tiwz7njGOpJblI75qunFxRb+bS4YjrEj8Pj8zD
M1bvr53otdeSkNVXkNQWbsixyhpKYBiRXIG6gOsdHSsoVUmyJoqRltFSqYhU3wEmIFKbpXaV9GXi
+9MWpvUN2gPMA/GrCYgD2Gf7Ht2o0QY+CZ3qzjWwL8X+o6kLKkvQLSWxg4K3FVyvbvteMSoJVqOK
u6iEaoGVqrlvIrRqsFVkfS/xB3zfY5a1FQ/MSr1kLhsDmqQQdXAho3ExmhCnCP5vlgFn/izGeZV0
bPFoeiRqLULxDjTr39nh6qJw6FxdL27c/wn0VfIjinGeW6uwG3/PFLh9A2Wa3AOyLnsw/T7PMusa
FytJqgFX5+7LhodbjcuC4ZZ2xWkQbiHOYzt1CiURC5ndfrg1lT9hJ0rcDMkh/+KPKFaBgg60el/8
bAS/a4ZodVnKhJNiUFK80xSiEiDv8uncKNr/OPIIT/XQB5+UpC8G/iU0+RwjQjklwAL0W6hZOSFj
1xw7Jc8ylvY+/hCzAG8mOkUPndcIdarLswOqTFV6XyDqDX4R7jYyAOrtJ8LNpJSMlduZ+KjfkTP8
UvwhSCxHRkJ0fRiRLqUqMtF38zKDVIJizQ1v9cDNm5jO5YDS0tBMHHxcoiSGgnhdfsbqTZl7PJlB
9phKW5VegqKdg9QiAhcfsQnYWOFrTLUYW5yVguzWKkLqNCg/jFCRDBrkcakPYKgtdAz5MrBzySjl
clk4y9TwZ3iBxAyL7lvIJazUFM9bAHKRBCOSepjMcehV7TivJJTRyBMlM2EnP4aBrqWbZomxMra7
RNFPZIxULqiDufZCbXxscNkCnOx76zCdVy+95bgxc2QLz8hqSjv0mHg5+yhT3w+soInsmd4DPdlo
dthV2Dby4R8NMmUD5eCBNTGzN4TZLN8VS+4vgNMeJ/5xT4Cj/GDPiGMN2m/C4gZx/TTc+wIMao4k
WH0SCmIwUEyoNYpWLujm+9e2vjlrKz/dLIMVNtcDagZbG2BZw5CWb8XGoPrpiwaf1i8vBDELqywg
kQ1gz5ArQlT9XNwv/vZC4nD5aSVCByP4tt2OiIzfDrcbM/T/yIKlA9luhHn+5sp7lIPnyMh7Jl8S
ZenJwfLnjAz193kAn5OW3msU4W8WVX4WtSz627dochHuzvvjmuoiSWpZ/uQHKr3M34q4iHJJiEUb
87GKRl+MdNyC1tHAQY0U7bcRsrSNSG1rG+FXMuupA8sfPjaX++gOyojj6KZMMebAHj/7PUlScaa5
TIQu0TTkY1NIEo+2LADnKgi2PmgO2FTh7fuYL8h4yEeJQJZVqE/dL8xW5lqtcanG0LKsc+kQ5duV
Ay1RVm7F3A+3DO71d7fskSADwL43o17cveXsvzz+jp4m4mh4UxZy/eSGmao/tnyQxRtjy4rF1W+6
MhaykPacIlox/t5zNL1EyCFAJ9pYlEhieJGE8mMWepj8f8B46Aehbz6jKshAryS50S/0pSkaMem0
TxYfsUG5zdDJk93BdXUN0ZIDlBaocF+uLFOQI+FAtaHowbluD1HU/DdK4YdrPKqscFWUewfKD7a8
GandH4lAyNh+rwW/Y0h+BAmzHAlJCjD1GuKwWkKrzvgX27DmbJVwjRNdM2TncJCf3LyXPQJYxcJA
KN+fIPCsReRcF+2NGLOlrRQzW7lZD6Tm3okGgHyVTNl4XYBdn3Rx4JJMqKKQu0klVzzXYKsITs+k
fFy2HxUZUrvBVVw8TVs3Ads8aQPFHcOME08xuK+OUgQG4ipxitfjn5ysao9pS3XsYBtun+oVx+1R
2YIGux4zhw4bXz0jh1wS8nuZnTz/nYtnn5HaQECMg5jV7nXp5iVvms7EWuIcQBLY4Z1CJW/O7Enj
FdJeAJ1WZPcucZwd2P4jK+csR/WrtBDopB/meB5lT0twEv9/zDpv0KX97CxVA6iyot21eSajO+CH
wPBTBsvJCEkgQY9cykdqQT5cBbZWi76T5/v572tPsOxa50aNDWZ/oB2XLRSXUNUAKJHcFfdFJ0/r
fXSouuiIbS+Euq8y374XnmRHY7rvt8SGlWaJp0hafsyWtdyZR5gIvm6sBf4PFblC4A0MEwWcdMet
Kv+W6iGwNxzaD2yOY7X18+R8E8TyWSyl4/yXMohc2FhGxfRN6Wd4JFOsJk34U/qAjT0585YYp3Qr
PQK/hf3kI5NsjtnUO4Y3DFZtPn1HOmy7cUg+HQWc9KQr9UF+8KwhMOd5c+m96a6RWYjEuuQqtsbv
CXLTt0ddahMl2YqL7ZtfS+HYYmWMFwzRryxgMWOiXc1xny1EZycDdUOcZqo8Skpi5gLeW0bdb3UU
Ta3S+wNdlh4tKIsT6NKUnaHZ3NkQ17bglQqNFNWjzafqmtdY74EfCHCcByeCeX0uAoWP4Hkg7JwB
QvUMVhDyf6K3LrfyvLtLtG589ULxe8TTZG/Sq2R+rfFM6YYh1wpnwnHpJYUj497h9sSRKicxaIzd
IePKmgZKFQGMExFHT+tzqaug990dvrpqOI1vWNgpT2ySSLjmdPEbvVyBmNK+qqT29zNPtjPYh7Bz
QWTpyyGfC0jGGcjIYjGrWJa5vkHevdlcGRFL3MPAwVgrkQJ4RB1HB20wEz8wsK+CZTfhQrVll+b1
+SCSokuwZSljzlG7nvlHfp1UwhNkNAaZI6HS+2Wpg8+8WLXuVoBdA+U+8Q0m+s2Rj0a+kfVNDcLo
cesiDbBX9Anr5Uw3y55lfgfO2M0UmehRnriep40RYiXc2KCYfWLl/pdhGApjC9JfV+3ILIE5LTGd
ZCRVxgQvG0wlFtXIVQQoLuVXnbPgthvHiCojWPWDwqxFmGNcn75Ma5m6TBeI60HpNQzxaoz0OVME
z9yc5TjDy4nt6NWHMv3BP20m37Euo4dX5T0I87OYqUIuR9+SIty4lScCCIquJly8YNQ5LioC5hQk
EPKG+taHL3yuhHpuSjSbc31F+e7p8DzUPcnP4LTHC16JmwInLeYJTLpNLANXUhTOWZsDP/EEgeIb
Nr0vvCsovSKcUZLmTCkt0B1QMjzwmEcHS+zB68TgwnIOzXgpUrHGBhJExd/tTs7HBmhsFb+kV5sK
+OpISmt3yQF+3KKJn/9IHNJDAXSmKu9jCGb2WmOVUE6/K/An3SoUUWZqYOoQXKQDDrva7rY9po3U
So3ux/iLi4IlkaRWnsO4Pg8+OmNTi3Y6HlB+gnvr7fJZ/YH+QLleo4VKCwrm1KPE4lt/Gg75utV0
of8APYS8C/jJwaKaytv9AkaT2YgIljfP0lqFCUVPBEFyat1EQUv6kW49CTco4tQfo9BuM6gAF/6c
iuHQL0BpRMHSEJ5KvT4XkJXQW4eIlIZH4PEr7MSFP2nLelTylFkxbnKu7KAVVHoUtty3sHic2tCy
z7GFhXSCUZcAaBe14nVUJvFLOdEZuZRYUSNUx6ZCRJ0MRYQrubHY/CMKbgvVUwSViRBXDzp+HwmF
ZhXiUpiWUvLzyNz04ZdMwoMITTqPDkpnVLg64YbA2CGHIcsFIb1xIcPOloNrUs7EpqCQuBVOoIHF
MltHfOAIoH5RtCf+oEe8Jm5uFw5erhd5F43srDG53jDfatBbbWXfeKcjvYz5VmbFOsmLZ2cSKmOi
83CPJ57mPng0VL9kWtnDadIgxEIgUwksJBUD+4K+ZUwa3jzk3LXFHftYSQihyfK6DHD2a8dxeUs6
yFGhIiQp4dL3XMHGB92g5fut/vv1CTQECKTGYVzqTHjmYTQKrwBGfcli72eYzQHJpupNM22s7O/3
ktVott+p6eyJmX2wIToqqZlD86SxBqlo1cESOXvYAHdB1W0S6pXjxvotKvjp1mC+UGv5HEMLQExm
DNLT7+0eKygy8z48mvDacH9nn319I0eLantRuOYXMqKYuoFPXdoaCP9RKi+qzGWR61u3UjgFzuzF
y5CHo46ttrW/tej3/kqTZnKC/bdiN9YM4SyqVyYJ/tq9TlMwN21K61ZqthAjKDdyYzsVM5HlN7f1
Lz83evu7lF7FEgovecpsoEQKahAYPMP95ZKh0xlZB4HG34RQOfg72e3IEhhMXJNxHp6fVPF6kDVY
EK01OrpoAzUL4XM9Iqd3ZEHsPkHv6pQ1ue1NmgppFbqg8AE/f5ubUxSdNxvCoLX7qROpFfpa+pWm
fpGE8vooi8nSnqi/FnTEBIY1WsEXQVzPYyl3cG2fwKuMBrL2Kb41kE17dCq5CqbM8RH0fByhOR74
8DIfJx1yxRtBiUzTGRM8r48aep58NVQy6QjG/8RtuR44J6XuAK+j3+aP7SWbyqyQj5WM91bA4HL+
HJEGmvkCBuJ8kcnGcH5OaS9MMNMVOOT9fY7h3b32jV0J0Db5ijX61YWRTCVTNXFAG8W5GDRU69Do
Ahvl5Gqg0ZSIKknXn0B4nnpXqV1NcvNyxlXEkCmYyr0/rI/zK0uU9HU/0vkS3qOqrYkPrPFZWUPh
gCw+3o+nX7q80N96K3X3S8Lq94ol9z6yQmlxwBj2Jhlryc6Aj4fYoJdozeg6N7OjpI9IZENtgH7P
Nzr4yrxKaN0pybSaqfdqwHlFL8cQGaeCJVrxL1faFJYeuxIliM264pD2mQzLl0tr9daKCjC6RRT4
GdjWYiENHB5Lp1MueqAxy+WOQi8zw9M+TWVdamgJ5iSyeYwKGRSQQglxWjS3ppIGZQQhb1tdp5Et
vlRKwlsdkueQGRociFRVK+iZ4VzzLnW9IQtleLiTaCX/f8OlTHrM5w8+Ccey9PZ8p76nFPjXD73m
fn62awmbC877k8Wy91EawuzzcKMMoqieun4DdwPNDT5jSLoJUjIT8X5NfB3ehk9IA8jIGl5GdR0t
eO6R0XBO4vF4SaLg4jWujfe+ItzRqMIi3Ev7FuSXgHevB/obL8wryOyl7QZ5JeIOHvyBG6W+Bn/F
xNd02w8J4nvJ4OADVK5iQlK3JgW7Ioc0QGQ2+h/8mo6PNsMpW5gyWngMWHdl6G7kk8njxb1EkRH7
0zuEZibsHicRs1iPL1Ci5u8YlGVVmYkcONSL2HIJOtjmW0YxF5Kf1PLYyGRZYVnKy8PKHZAuGXSP
870n0IIhPb2EGuF0vwIaXzk0kl3qO9uELkGJSaCf3B/0EV8UfbpLwPGcl/3lBfvXPFh+uktCiCig
n8rkBnRo0mUmqMa6TbB7/8VWXgJ1lMieg1RNL21xHHhnMdkWIlU526v908liCa/TBJyxjaV2EXvs
qg54w52JOHmzlQGwW7HnpFOTI4Kth2EsJaX2o3lWahTvjp4X2vf/4fgH4/rnR1wQjRE+hVtQvGKS
6ZI2sqABj/VsIsEsjVrysm80GNjEsM+1r45LM8w+cO56UgJAyFyuqVjlY1mqCNN2mNn4e9OAjIpk
3U4SXB+jO3+f+mVkMPMvI6RZzjT+8D9JJEf98SeGv4GhVxYV8t73G3uXQrS0n6qGwSrXnpOmC2BL
eeSEdg36X3vDW4zWR3HENicJ1pT0vMamRRyxJPvAnmwZ7K60kbaNynns443hKc/VS127oFZmpD9l
R2KXi9BpUofdYIr+wdbi3R8cucLQ4/2xkZxlodxzxSZ/SvKrcFwrXfwAHCRrgSpGdLqFGkPxPzq0
qpRrWg06rmj5dBde1MgRHcfqQx8k/5BvMiZh+WkASWIwbYQPL186HCZ5gcIl3PGNO3YdOpboJ1Uc
3pFh2dBd8uGWEmi7yFm6NfBE2mV+BXcJfO2/pFY1duBdwB5GhElNN0MZz45qfRTSMiRyIk/m/yp/
AyEvVn7mLrJ62fejMpWxwxSpEr5UwyLBidOnenbUEU+5c3BQyffR2gtfchllvEN+EksA+6lU3zqL
6aSVVj9t73T/BFmJlfp72pvNapJAYcihDe6ALifSYQLYtEpqRAYpg5iGRleKods+ug8RbdOqONv6
VUqaX/S9XjSfMXdcsviANnHeP2g0T2ZoZuCznpiBQMJiSC52Zdf6/E/z5DTB22iLwiBCPb+MeXsH
xM89aVSqhcRLEg4CMSUvrVEoum03S8oc/5c8GGHQGhTeICPiecZSbzEfD4kWLP0tjHXgtm4r2WLn
tfhC/hVS3bxiTkNjxZAJHvtMPoWcyNyxIphQ8j61BK1fDZqKFLSM2GlBCg85sYO30AYabvil5ab2
pHJg+bqZdK7siL181DZ+/aef7pRv5A5CvQ8hHINDEZcMHM9bbXaTcGW/Uz7bYZREzzvtgKjvX4Jo
YI72mG3oojE6aggpHf+P+mOSWVWU/iy25Ac8B34xxoQaaTOBdKVeBs9/AppSymzd8Ii54juYVxMg
piG2SVYiuX/UqFFzUqVUtiAT9sTzPVVTiWrfcKHUAyJXlHPcH8M+mEN95MiC4ik3FRXkzirV9srn
PhsdDR7TeQxXSywYceQ0Vq5O+JAajinwQ0V9AGPA+b6AlTe+xJs6YOK0lx0ICPYj3mGyFBMdJPW2
zNnFs0goS46ahqY44wrCxz08atY3s0OVcF4Xge3BMYSChoAh/LNVPm9SAMQuTEc4z3IG2MdZpXWA
D3Eu7fvm7pYOWEQ1tOzv1XcTEq9ibWsS16Yskt03oNb7KZCdufRK8I4HWvJ0PmIsS5dRx62ZZ/UL
hBbDS2nY2qmMhy/2fM3Cdc3KxrqOQfqL3EUbQhYtk4Oyzi37mRPHQiJYi6PRzLBss5+1eH3cubrQ
jbDec/4jjnOkomuuWglfCmEG/f/ykC4J1h6C9Ug6RiRJjGFTinP982n4ojOW9CRWS9aFtxIcE9E+
ZJruJJXOV8AEVw8d1JzCrij0mdi51Ar7RZM+PMvdbdLEBGiODYhJeSjJdYvfk/VScBziVix5cGXw
6WQCSfAXSowQl/lk4VKH3gPDArlHf6iyEdTn4sLxs55WQ/zYtKtyRIq/n4D2iKXOv4Vfgdz0eTQ3
8ZeQTCO/5rJfG+44oJ821Eqsu7cE8mR+7cPICJSfut4l9lFPWXMhvsDT6miaVJqQdleJBlCf9/iA
7INgPotqoqM1WygavmF/cb3wEtRKIMZMX/XbQQE5UtLAfZjj5ePYpaWP5H9U97ToWA+IH0GSyNrA
KyUgFGA8HSUi3bhKryzLykgxdzUOnxrjTzvDoxTD5LrLzB/UqkzTW7dRt7dmxIkc6MIyIo7h35gc
DhEOO9ec3oC7p6T7S4/GJ0mXLdTtehxQ0AuaS8Yb42PZS5+1Ql6Db2QYU6vqWujC7HKUf9KnvJx0
Rjl0rR2O+niwEoU3v4OZPF553ewLbTU2/q6F28Tm6wB3p61swJviFF0ry96HAfrELZjaPOheP+Qn
zGbyAc3h15ikRxU8+qK582BC8lZc9NhGDlvwZD1s8BMHC7YZP0YrEEjvSiV01nDiv8qMLzY0Q93E
5kajwNog8DSttDSipZ0dYHAIrH0fsWB3VrwZwCUd1jP0U9iuDF6ZobONN+d0eXQrm1knePsC8QtB
t03xCUMVe/CntTFjRYnWUkh5oz1uXUgLqkaQtxUdDkHF3dNHJ+UhsclVlfOjh+K9qQ7LEq47gZfD
a7OPJo8dcfNs2qEPnYBV+N6f5wvJhMtzLuVxwmmELoh4rmRYvU5RL1GqymOPtI8osx3SY8rprGbE
SlM9V3VARSfs3AR/hTi6thaLaLcM7jsfCFIZXQOkk/kVejG7OuDA8GdtFeacFz9UxCbYheQEAAlu
KcGwpw2tYClwz6knRe6h39zWgoKWnfoRnml6Os6ax37rShjRIwyghB10RFzSiTXSgQAycdW4v5jl
SCuK2TxUEkgAi0jGpIFT7+X/zInrUZ9OCFv/qmlXlJhKNYv7zdqeZ7lXCqeq2S/Bznq6lmDUJRsG
8DC34sqgblIi6P8FdBSalBHSUc/oUN/fde+MGb/c3yomTdhCSpp1GPczrumT+bUkPlWoRETJk5UH
RsRKloEdjkgg0qs+HNIuEcLP7wuNghYD6kRb1E7A5PYI9yk8INP4Y7FsgZE7PuGec9uUvV5QgRGL
sfFe9IVSw2F2Z363QPUatv1hHt0VjZBGrDRoCk8xGzNtJGm+tr7ebPGLedKS0d+gatE2zdswMfJI
TDl0a5UkV2n35f0+pgYr2mSkRZBWzZrFkOLbwHTvoWhkO5a4QaUyNDTCyTwxObD41yhdq57b3S5h
gB+2FyG4dGC2rBvVrtwAaK9q4RMw6+NKPUn0j/kW+Bjt1tl5P2g3/l2Byv/TaMaIx99IF65AnKp4
ypYkMqbNiXXdlpppZz+gTCU9CULXXwZWaLyHV4F/d2B65hFE6LZmiu5AdM5SKRcrsT/SX7YCiL2B
eNp6GZtmA5UFvK4MPpMAI9LSloxwlxSh/bRhyeIHWJI3Ctb8kKRp1yi2nEXz521nri6nn64hUxOC
0Y2Yh3+tIcY7vKQDQxZeJI7WztOKXv9BeQplwzND/hlTi5OT05uVvE9G3GJfMraRn3WFd8rCVe9R
lZAnCwo+dh+vH+6ybSa5/YK82kXNKpZPLfK3oRLqSKFv0BhO9kKpHUzHSrRwHVCra1ig6RAceobj
jBNlm06PoLb10YHrzHwe6v1VnsjADbJTXPQPt8VGvJN3xeUdnf460KcS+FAmaetYAt5lgiW7kvRC
kXRgwa9zznpE98tCExCKYsC1kpBPPiWAbQrChY9f/YHVDO1NNrj0ePoJ7hWr8y7MK69rpMOUopWp
E7WUL1qhSXFzdn+6xUh3zeQ2q9qLJBD0eI3SrKmyBlhZfhfC5fi4+4YQgYV5c6TI/gELjpMNbm/h
SruvKVwV8/Qt4nwGu7YbYywG/gAO/loAdrDarVtZkOXiob+mzudrNgFyH6myNBofeEbz0hMHzRCZ
YNtsGKr7Ld2Vhk/FdDM0inPKBk+i/2rcPVRSjoQV8bLmIaiB8AfDgZee0SGwCJKPjgbDg9WEla05
K1FQMF0afY7SVqjZOIL0ZJgjEFEi2axKYLAyIThqUpiaM23GD/qfQIdG/q2/JWV9Bue8+rIsw7vu
nr6Ovejctbm5vF2utZ2Owcs/shT5ba18hLgayOxxYqDGAFj0nRRPxk00Q2VtY4nN59moah78/FJi
7xtzFOCzCe1AjQrkrY7Iuw0qIM0YSy4zEwzVQB+7dBrsXXyK3Hqn84PVafLozCaSSJP/wpPE0zXv
Knrmh8o4pjVRlQWplmEgf+Tbz+JAqoD+peVvhquOKC9DnChMRyvHhTIDESQ9Fgmw9otWA/dcX1Mm
M1NLZEFRBb/mahCfH+58IRk7zuIfc44UXM05LUU5t0eg7oheWc16lkXNa1F3oOQRDYnDEaIl66Ln
mXdzkEFga/RaaOKbvX+3Z2tNQkLT0pgPikzKhhBc9txMQ8Ic5Rcg+vBQ5HT0vPAgMf80Ub3aDv3q
+fLQRO7C77mrXdAi/1wLeAIKNd/30Y8wbh391yCgooBlH7U5zvsQZV7+zaNZgfMpqCoouyJxLI/+
79lmBcGkwHUhUUFso9npj4g7gtAoEIFX52HV18hBS8u8kL0hf9NIwMaLs0p3qqb9raQLyyetyERV
1hK/wjBztkgjjmTt8yGHvU1l0C3Zt3LFhvn2or9FWUrfTr+5KX7JNUEuA+ZcccHGUqGayAhybcef
cHwyoh/KJWb+e3vNeATlkb4WiQplycMhEOijcgho/A39VyvD3cMpKj2JCLAkZva7S6oVT50SPz51
SfXybvWJgt1YzHtZ1zT9eWvgRG+SbXJcdPKerexw3PHM5YQi9jpDNmQ7g53RL/FCksAs4/wO4SQI
cjR9NVbbO6ntA4guPGtrF/H0wu78omRZjWdblQwG13KFNJrBpPo0E59p2yJgyN2t7THy0Xs6StxJ
pZ5ZvlWe3+4ZLG26tkgfF6VUkqwmmjEFBk0byYDWHnQ0qiq7J3VGtauNA8wropnqM/3fTBZz9M36
CG1swaCoP4LMHqVamjMokrSerh1OQl0ARNrh7X/B6StjWEq6eeKOfJnmwritlqTs0wEsIix0kyDz
qQXPofXkKpgq7t4CuBaEMK56rGlJNrzDph/EtO1ILzM0LyWrrB4lhlUM64m9X6MP70qato0NB4gN
1h/RzQn0GjQbGyIG968IsiICiFSW3LVKVU82T4WIa5nCiyuqqSXEw9mwgR+j1qPEevnsg+8DRpye
w3tF2jilhrEJGcUesOtiF2sfBszrzjXT8NS5/wVn8Ck+Sk1eZtV/DoaX0OghUwmplfx7w6z2wRfy
OXuKa+KimxGSqxMeFwMSovFoUjuYIeh2MJBDdV+OPdcYsfxsPNhqtaiRNaYGxRfoEhN9yQlVev6/
ryJCvNQCVi3fd/sb0MobacMoGQ4pC2yMvxMQXnLpR+XDHQnF5rBBKWs1Bs5Cp3ERlZ2Gz7wRYGyE
Xt9K7B9FXGs9Z4Oo2Jsu3lgL4dswQ66Lh3yjbI7R2+40AWMvGKXLA6YWdRLe79pzFiul3M+GLbBi
jvSTsyIp5a4JGx9eZUOpR4AkzMjWb8h8eJ+ErvYbnrl37ilQFQrvhzCHVhCTEtDg2YfJQRwiVIO2
uZSuhB6mT8bFWehObWZQqSjwXTspJKf96/Jmdxr5WWa1Vb9KdTtRzDnBQc1jlCypDz4mP0/PoWCu
EKqypur7eslM+OonFwNyYgnaBypj9LWeP9fZe58xgTiqFbcuamrZxTXDAMEm3uap1ZcJr0wGVc+G
8XMEk6Q6P8fw6R46XLTPiY6RYLv2NGsFpC3bJpyn5wqbpb1YL9PlXTBa80O4KMG/pc7Wb0/+iifq
ZWcxTATTNYTHHZ/ZE+kT+7ZJQoex0506lHceBzFdBZX2rCW1IGvvdS9yJDy7qUgT+dz/Q6RkX5g5
f0Mzjq7AU+wbTDVf1p9T9rG8EU5roK6gwGjedchLjEB3crvR+eL0GPhN78MkBV9V481JTK8ql6eM
4XDBHZb2AO0Ym7q4I9BkXx5wyr/8UK0TJEAowIOEmyLSie7004odAsVNL8LgUSK0KTNsn7Zxdidp
OKA32mgWtPkza1DND3f9EiK1uUo6dwksvaTDEZh9ApdxaLfKhsb0JnceKsOx5myEjt1/MdYow5LR
BCQmVtu7X0CgJsG58TIFEJ2R0rArxIZHEqrcDvENNkzoPQ/bc0YS0HUelTEVpA4MjRDTSH1VIZRQ
ueJ4Gbr+AmMLsmyApbGjp92y7ROYJGNFg4m/X6nrv7VKMPwNzkFg9mx6f0yL62WNC5tjqxBcd1iN
HM/9XqV3+NChcK5UP+S48eDuqzpBl3Rw8YCApfw7cvdQer6MUha3rHBIx4Gd+l0SmMBvP3qPpkRu
EfjrtAztJ3+Hrsx1dIEnuIId9+TCTO9ve+L0VYU2lz3fiQ4Y/2uQKDg49q5nCtUABssNu5NbQNOj
qPxLzQEgnNG8viznhZ/3yQZdpX1Sj2A4SzXexFHTcdlMCwu9bvANidVMK8gKZdNmZCskflLNfoIv
gW/as5ygyoDEnxl48NVciIRbM34wPaIDO7LDinSC7kDeKDPNHUMS5phUJSqql0TizP23eBIDA33V
vSZhqPC+z4xZH5S55UVDRijB6T0+IBVBeOroW13Yf7MQ4+Be5VdE78gBQfKJ6H6sTrCgIzCMb/1m
oeXDvjcYbyJ+r/6pl0guaeL86+URQCEkQ6GbmINwI3mWY4zxjAB9bcCutCyKSFrJNfAhRud/ht+f
Gy6PKTTvXZNp2UEFNHUidITkoy9aHL7Q0RCmTzPkunBOMSzdidtdPqRVgwvRpb7Krvms2ZKjX4aQ
qeAXW0V+k84Dsg16Tf+iO/K3hIeCN6XSc8MElVI+Y4rkZKoWnMtH8FUs0nJnyAyQsvUanF+Y4jy0
TG9HVHuyBV+zULDNDQit8Ow8/xr4OvU3W4CsKoePxDMgQLTEDaixnC3jXag95Xh1sn0/qkJmSU5n
ahMqVyf05GWEtGdAWMykxgURuITL80hErI81exBYL07mrWq/WtQkbVj00ip5VLD/X0iBG4gMwMXD
TmrKMr90yHHoJj0GgFbQeJ+ypsWPe+0E2SToG5FhiIiqHJFTfT6YYci2vt7AlNbzDFfjQc9Sx7RW
ffjQa64S49ApTToVUI2FQs6dUPysqlt2N86WmLUajGiGvqyIE/OmfOM6f+o7D/KG5hhsYOqT2yD5
bkyrhsyIMyHlQiNccdgV3KlI6k2ZzNCu2NkrC8MFnhPpsY3e8gF+ihkPXCNXEW5NJoKwfiMYN8Sg
ZWugezzjvb462trOUNVljUMSPN4SPV8wHuxfzvfb5mwjWmSR4gYF3ECLcUi/O1FMujlFDjetm+HJ
yym+u8CLYttRkFHtqu6ozxuQVt8CRoMYbQEilGRGNTWVCiOBH6qa4f468TebARucIBB/5FMYfC5Z
Mul1Ll2zukokfF9kDae1EwNBFMzxV/94V8SotoYrOe5x+r4feXTTBJm2uWk0u4pVe6rD0zasPKor
QQfZGpctQtXDDFQXtbt+5ICahtS0OEMjtZ8f1Gvo+0QtSkYxsn1JvS5Q68N1Auh59oA+iO+GnxBA
nTuZu+j/ZGZqlW+DL23i3OFrkIZwIWOj4lbdtpzL6b7kINdQYN5hAUdpNu1hATkfvvdON45IjUUX
LwfAcJ932jNKzPxUyI9M7YRctaRgGI7pQpViKTzyyOi+qZBblCHmWdAZFND7QRKxJHGk3dOp5P7v
yLqhdy6GViKXIfLUizlAKJCydlcxenpDRNXFEUOGHyNrSiYeU3KAfVDtj+FVe8DnkpvLbANq+rH5
1h082/7nCjwwncUQvLFnOqdjvhMXETU7sSyXuNA8GuMi5D9h1GQhGzrZHhBvUA+2Jcqyk6H3YBLk
jVzhU0yPE3zxSlhy1mNFEDrbDuODhX0icUUx4pIn1uQdrDDsKCjccJ6djZfWYSErbUV/i0SPXvOz
JZDO4RUXEEK+UAM+vtr1xnG1plULoKXroH7zpuC+ygYkXjMsCBqOTIDDYT/yrYnODQ1xiFS/T6RS
x+K+Yg76DNIVPnHa+L4BhyL2d1oukDh/kUheu2ZSDCrKsrG98e/XBcxhV951DmG6su35sO3jr6Op
dJ6sa3UWid/MqinaIaGvmMuopuSLdtzyCIJExDyrbX/NvhweMZqyNq1JSjYfA9o5d47BwPfJ4Hmb
M5rTbT46zr6Amx1iZixrh9uEo6lz8CbiF0YkA7fw0QmD7AjvSl+fxsHw5BQZsfmFNCArpaqWpNtr
zIRRsuSR8x+iUFD9IQPC+kp98lPkeXuBo42K3RwPA8XVfhumNti2bBC7Jp0h02UEw1eSkez+UOfF
xh8MpBigpjJ6lN7a25HtU4Cn7+5rvA/3gURwVeL8nuUnrxt/99uYmq8fJWw8Fv16TyFsczSQWnmC
6hXmQ2BSeVS+hX6BJnVpDyglv8pf9XPbAYHp77zrUsfFGJf1l6SfuLzBPLXTKFINXNoSISegx7Lu
gsO8BD+CZLnDMlnx0h0DDlL2wVX4ebYcr6RoaoRj8Kv/2fmcyt5huqo+WYtkCfZ3SiaI6qWFndmN
oyY+a6amMqbWKxb/i94fjupZaVnZQzN7dORJccomjWwP1JkHd6g5MVk0k9ELL+T1Om7OAVngkbur
I4iCmMWagfAKfj9RkxOLGOkzQWt0xvYJ1RE6xsUYckVRD4g8ewFpwaG1KT38Dj7cwYd8hVb8Oh+2
bYPAPlTMFZgGhJsSlaUXc6oteOr69rill2vitD8rTURBzzkbEn1sWyFhG6ErbNogM7rhR8TV93nT
tHXfxUdeEiucZ512qR/KBIG0v/5ZPLnbQdjjLUTDYlvUFgOgzGsXNPN863Q4yO5WJleJHpdLLA8k
xzfKX3qyCNGc+cQm6I31cQWDjeB9ZP8UuBWPlrCyqJ1HGZ/PYwtOY1cMpuF1UPvYDiOAA0uyrxnu
vgZDSwjMEVZWszi1QyMXs/SxoJjn493TARWaLBuZZOtXb6MDJgvE7fvNTLpdiA4wYRcDrMnl0PM0
+I4M0f89VO+TQlUnsiIEBkiv0n1ikZDgCkwk8zYyEeW9zgz/DqQLDiXdW6x2BswuuIKDdC/X1YqU
mDZ2GYuqI/Ly565um72r6KBMo1OkhKkOG/X9OtS8i3vZkQX4jXef+3CozFHNeLKdshmSNmpObn6z
W6kWAmYu9GD/d3kfeR5maUj3IAxHbjDj1/Lv02zaDwqtvX5xpgU0m3tpAQ5ZtD2Fxt+vOXNzovUZ
IQl8OZmQ5yd1safS5sNXhDGmXHEPcsJ+WmmV1XEQcIn0DTvee3qwTchfn2+XvM8zkpI7cwGACs5S
gEe9eSZeRmaYrz7NhtIBz0BWvmcK5CSLntXDBBcid6NmtdTXAcDxNa12V7Bd5K6F8Y9x7ui/zsoC
92s/IfsvK1/XRTPI3/KL07GU/99GeQDTZ7+Fw7hlsqcRkmHa8p/7nzHD7J25fyy5wfpkVuffVEso
JTEz2rBlGjJ9CWjxe1N9hpPGFv4wGTIVyJrq2ObxCwyVw4RCxuFjm6PetU69iUHOnQjiY92eqNiw
OnrP1INRXdR+5xuJ8g4c511fCKdzapPzQCxb0+qlJ1deu755qiqzh0w0cjaeSdSI4MVeEw/eXRqm
SbtE+chkVHxj8bJU/16q7IbKqTxRt1v6zuX75dy51EocRmijvmkZSXxRyVmQZ7ixCSdf2o5F8rxb
LhrI2VrG/uOS6w/6F8Pj2+C9RU9+xe6vebPoo4uK1QJdSMYk39nQ8bfZT18X1JXVVXJGsiZCJLVJ
ju55Cci/OlyYj4OHNIi2qxJ3soubUEVcL/zS6QkauDoPfygBBKHugotd64Nw3RZkiu/F609Wphjr
AhHkm+DNJNGyMfaQwr0bPGTMIPAV2rMgI73O1IigIedvS5PSZiiHBGBP2NSn92MuWC/Y159+WCu4
4gaj22Tys5I/y5qLi5r2bMzsmPodtjRQ/a0VW1PSnsqCMAGwhtnz/TcowqFAQ5o+alkPnBcl3Fq+
weYKjlTlVyqe7g58cSmggvj4oPMICd3ftBrRC1+yI8Spb1u6fVhTZcpy8VjMDxlKUYL6HWXPzbwF
UK8UHJD9SDaS2oj9rigfVrBFkWfEVUSJ25AkITGJJMDhM93urZCz5l0xdM4/HoVLWeK8ltXqygCE
I0FPoveGpMNhIL81aqa2lLblcbiZrhoSOAI588uoq0kghQUR1ARAo8txtaByNiZ/vL5fK1znZ2IQ
T09RlctbDO7zD7gAtERRYNJAqVJwpPasoRwJWiJWlmcbGwG94HfKS2foSIZ0Qc7SfzRH7uuJ8prP
/t3rG5pTEliagEEygD/PZIAjuoDlDeSIF474bein5ojMo9clxvAt62Ey9RkWT1lYVA0pKqRRGRno
V15rxm0Zjr2J3fLz4DCjSXakBrA6tHZKuwYvotMh8wAjkKo998ooPisVpJazHsF0GAKKJb5Y/vr9
3bHzjAcAwLPPfuoddiGPrdY8BOjr01n6PqSXS8BT1bL7dkpg+PMtpGiJJXaoMnWZvLRkHd6rezZL
HPtEsVi32i1nttF8MAWGDeRr5Qw+ceNW4u+XifGlRzuXKYhSIihWaTpgZE5IR4f0ycRwysGBejNF
wAxOwUGTqJ2ZQw145dHBPokvk+Gn3mC016gTqEDX9+rIb5XDlnjENVKI3gJJM5tw4qpceQk6eGwZ
Iva6g2D3nWMEepWa5GiDaaTmBPNw9FaOTYh4MreuNNuR8BP75xHwkc5SP8HBUC2dCNxIlWB7nJIY
AIVxVjwVFG4xote5qDAI7cEonWS8jhm2MFOx9GJX2j+qMKQ5SFlExWkSI+G0b/LkMJ38wDUCQgPW
cXO84mWsAFjR0uHOuNWDicv3fApYN05nRD2mdNyOqFPjcSxJ8fBnzXepdDk2WF1kB+3K5M5WMA+h
7EMAxoeCOjT4+4B8X4pZ9sSsiFP08gLP7ZHcvL4ngz/31cod9x9CuuPWYNVxDl2BAH20q/n+IVrW
d+a4sCNkOMlAFAd9gG9ri27rYTorAHZtkEfEkqGJOSSu2ShoGO0+VLsD8cR7a6XhK24iLJFjTpIf
j1ih0+yLSeSsAOcbEIs2AfN5ACB6Oxp/uFU3yuWUNQgXpN52Tezl+UONL1MpVYW2vbD+lwcYlLGW
IF6nb57zP9CefcFakPKbLH2l1YCHIogeASln0ME+qMwACxRbDbqPc6U64kTmPZ7Aec1WOvzgpEqT
ILI8QdKQCS0vj8P4kem6N/g5VtfbdC86CO/e60+Fwjs6Dbaa13ppYgOzdeAe8LAZ5WtiUkIXn7lF
E452iBWlR8PYa9/NXqcdep8dHrdOWzfH3joF5QGULdzbqFM1UYRRx+WKdDVG7WGsiR47sF1jWWq6
kUNWvw8sMZ6zEa7ZKgg2JqVwle74YAPUIlNNx3Q0FV7ErfTa2FE9O5KskuxRoijLR8YoaMBkz4pC
duzduGtAQA/q8a0R23wZ4U0n+S/EteKhOIejiZCLUELt5Du0lP3C9crOAQGbLhTY+ztv/9iGO10U
MRGaZFDtWLhx/hx6w9JNbPT8OML2OrJH4wcx/+59ojNgDFX5xnKs1YUc2Sp/xn9Mv6UFgrASTRUo
GIPGiwBpPpDF1orxTWA3gbuThrO/9KVtPv+jhcdxuFoq6P0s7d8NPj1O2WEdpMI/EnYtp41oF04A
X9WcgbTRy7O7B3r0TaapgBLjBcx1wXWkSsIRpKmHdwSQo+b0TWhutmDCrSR1ktzVkJF7aiE21ZFs
MrnypD65yHtovg5j4tCRWmEo/p7DVhf4eqZSAwU7XQCm0QIKIf++A070kTfc4nuzCcZevDkU/ki4
a4AkSyAAGBinC63pWJj8WIpAtKOSvXRs9u6lr7Jy+H87GJDviswSHu4F1eiOyEDayPt6pzuAGcSL
qYZoto4S1ca/TukEKiLlavMp4S9SyZAguOtk5WQxBsMyJQxBz5TZHyYiqG0VpslBIclIj/Ibm7yn
yfd4WhJdZ4vou0aA2s/kkuc6CxcmTVFWq7MPtU7pcvNBQi6GcIUL147gMmaPB+fF9iGWv8iS5qMt
aK9wbLq/e+7P3lnTFRH21TQft7IXquqVmPoYwseeNPwtC06mBcJG7vidSntznKDZAMxzE15wlv9Q
takiE6FaBJLy2UsairmaAA7i0L0FqweM7MBPjRI0/Mue33w8BoPU5TeJxjuKiv8OSvFxezcuWesr
59Db2ONK5H5bbF1UBpny1F8GIuT250PTbuT5ypSVmpDT8EP34QX5v/knSsXpq8r84YK1tuZfxl2C
DJR5ot5JZ44w59th4ANhq16/S35VkjMXhPDzlIl5QzfgGy1zkTIgm6ixZxpPKmtArCuAW2d78Gxy
86kPTNwuZDFZ3xznOA/sdkdDRJjpLJpIFI72EJwTMxDcLOe/1FwCnY9K5a6HpbXyaRyg6duMZYed
Sj/hUzq0Cy2SRlsOl7t1xMpTBtNi6FOSMg8jB3cn2zs5gh0rlnBeinOA034KsjyUadZZUGth8Kt4
+oqA3T+rM0szFCz7C2oodPn16NZnr7dRr+Lc1FRclCp6rthveGrv6pw/31X1j95SlUb+asY1i6Ez
55MOnq8GkxAb4EekYKdUwSKQcLvAuebdrLVvchRVgovwnl6Cj+9SKXv7BDs2wory3cEL47ci64gd
K94s9vbgvmRzo3PF4yqJlJkNjxzlWaCKHLuf6YgzPcRj30Z9KOABQz2NB2xQfaiSti+RLgM+s6b7
ALyAo7rpC07CbVW/3XfSXpR+AaLr7RoP3rnuAsqizAx6u5tqLAQA+ZJNIXtrI3GlTwO/GPoa6N1m
qCRZNYDUuoGiJI+SEcYa6+9xRxdNkCnl8QWOzi7X4IIr10q96GtsURffjUPqTkrSGlowdtP72p+W
n+WWnH09CJE0z5cMQwoDqBWiGbBmuCNQISIwJnNnovVIeUht6bMTlBx97XF3ZpjJebX5nb7fY40J
+eZg/7f0FiRm/LzGK2u+TB9244LkfKVmR+83HRMeTDOg4YN/snuIXJWyW2eJkCr3ISjYayIxL3g0
RxRbFzaHps1HF8qXvJ4sHs4QRjwJriGd5bXMiqs/kpuD2Wu6sSR7LzOOjEbJp549UHkrz7B8lGNP
AzUZ5FKxu7ghnlmawou+PSj6SkD2awKZhjmxAwGO5S7F133GNeMnZKuAZnGjb7kJ8QztJ3cZt/WN
EoVYn+ks2/tswhZJxM14Z30U7x9IHP2TQkN6NEErSMZRsy4trc5Y9lqviG1WFINCwG6kk2ENIoAf
L/g45Bld5vy95S6RNpEK5NSZ25jnLeeZZn3gEbqS7pfn2qtVfjYNm4ViHhvzCzgmoJeFsQ36HLwJ
LP0MGypMoAUMhQzM6pbjLuMATUlEmptuzLtBD7GPIb6OSrmRS0zSqbtE/tprAtenfWM+mIGHGmaV
4/uZl8p90U4ITYNJBOynmfyrKeDym+nD2Pz7QFsiWCDcnOBcpOdGmb0Q+R08slyVneajdL5xpNir
j/JjbH0NHCsL0h7y1g+GTolX2JLOwZIfmmu8DtPxnTcMbqFpqiB3kXpzRZluK9SvCuBEfG4p6xb8
71xV2kVA1FzyAkj+37WUTThiO0bhdRNe7TTgeo2m3scfjNecuyNfSQvBWvGGhOjwaDpAj1X1RQLR
xVRUXPrU6P5K80SHoDJ4oT9C3MjJOhlYQ0aZUUa6fZJ7FRLw6fna+XVkVlxGeYkkDB2NlMOtM3E0
It12OU5aRu0mXXi4KYruLZU3qjFwreS8urhfYAfEsxU0IEPuZzmDU0j7neJlCuVoKX5us8OXy37Y
VI3ClbozalgupPTZqsoobcU8StFHClp363hTvp2eJpUu1JbyIVFlwQ5QPySzwGmERoPkthST/W1E
XfcHiDxtcNYlv9dgynKxjWlmTbn06zC3NrMCFKIzQeo/NVzwO9aJsez6bF4ntNW0bbvwPyyG0wX/
ZyNOhh63UF1MDtWc2EyeKNZIMbBOpqJDcdywGi9TWUMhitloyT84l7skjM8Q6Obsn3u5wsXwTuB/
JV4+paY/6hL686iD1pe9zZ+J6m4681CApdyNdhkOL0yUP9qoGPVCeSArsg/54ppTmYRyhER6Jfxx
+HSV5JlZOAIMuU3sZLxr4Quvfj6IVygWdcfkaZr9pkf2PoSSrOZNMult2IcoMjtPtEkoWRFej7Dk
9pLMGHBSH2A83aWl2dhD1eBmsGb2bYZ9Y8eU+sUOYzqNgxWuEniOyNHic1LhvUbTQ3MjHRsbsfvS
BeoHxAtRaHAMsU8k6bvVgjJ7dxzvbHt6Pk8Tp0keNoCPTI6HYwdBSs/swVo6eWmM572cClMv1tPo
qxcgq0pUZmSwOp+Ru8uC34UnwLwoOlkMhUlQH3YU4L1ljlI5BiZJ6mg4oOrTkfh4zi+laxKie3sd
2edE8BagkuAr9Ju7Lmm5qhNUNLoF1wE7/kSG34aJWc1KLxnfnFYb0ik6y8IXHZDEyVxrkIbN399T
wW97Vmuke61LPkyf5voWlTIiSowV4XXMK9+SV1lGehw25r2lZtK3tmobzmz7gR0+8X/uO2QJ5vYn
yJqHfCGeMnoEfVSW8jyCqcAvckfy4vUYngtudSLUiF2asUY3ySkvYIpdGxvfRPaUOV9wJrT56k0i
oR7U0A8ObTtXdqRwi3P+ME4R8Plob1mir93wOedexY9fmB8RqN8YwqtWtZOROQEv29ffTirc2dWD
MPBm87DMFiNLrldm8gaH/Auv3LZt9dDIIXt8eNZ3SRIzWsij1MQVkGsyHEkOI3oIzzCW4DqfDVYl
F7z3//N6I3wGyjv/N9bsZPHEVtKHKrtAUJ/UOlXyh6LOwjQpPQCws1iV662wHCysIJNaAaSFD1R3
PtuXxCrfGuA1uZtWAdEMX8xCELp2ANh1HV/TcdLpbgXu5dTlDLFqPDkuS/bUO7ZOt2GEMhEcut3P
CWdZzp67cRQVxPo+CkJrAIjkBETP4utDGWKDz5LHTx86PObqoddgtB7kH97o1IsBTQm50reJPxEi
TqFregPMiJ1tlVMBuGabIOp7jhoKF8uIHMJbwriC6IaNdu1tYclmiY+KGhsJ95eZcnuMF4X+VsBo
ntbgas9yBC5Zx4HWr5BwX09lrMvnc9BxVf9Z/ONZm1O9i0xZ5lxQ3Sfly3nQoJGHRhiu/z2pngho
8XH4SXq0VRfPXDD5vlare1w7Eei2OBkYuVvp14fzcbSJDOcsrTlicfKUTdpiC9v9r4iYW1EKFivg
TCIe2FZ9YIEwwi1xhvljMjyL4jZlPwPXo6CgSOIx4YFMdsddnM3RT5GeYHFZW+9MssmweLcqUAa6
B5jAXfzdzWvCiKKrM4gNEwHFk/NRpZrgRXbl07nzXXP+mlV4SSp7FMO2hgwoGyz890rhmz7b3U7l
Q2M56lHgwU/CZAYky9834zkzhfi00RvRrxLOC+jdG11Fu8AEoZ2Li00FEtn92HkyS+z0b8GPabTY
coXSTOrb5TDfFpTAHWL6RP5VH76ULywS+AQ9TaPb76fvaCfOXudjd+gQH/VQuR7Rb2+BYaUO7igh
2+OgvGaVfidHn4+wIvCcukkwgI8Nh9it/Ji+ivWrCvvB5wSeXu+PSD/61/eYUo35xbOTnW2i+OcO
ejz0FVatwqzhGDJnmMl6T6CZ9UNFHPVMJhj2C+Fu+W+80MqIu4CyxaA2V0RZKnUxysEPQ+hc47VI
/QkXA/t76pd6DWi0KVYspx4FxXM3Zpin4OQiVV+Xr78wlqUek2gvJ6FdpwdXas1VP/DSBZC6Vy0k
UKLtBEayAFeKlU0kUux+QquEYc82Lle1s2ryZIJkF9pcdaR0LnFP/Gy3RKNHSIfWWDJZrOu9lKBu
ez1ghkthDbWKGok4+VFEmD4JKWg3ASYq2244M31aDOUTtLs0rOenBT5hg46K2yxp3PB8Go9204Ty
Fkhrkqt7hdy9saWW5X0bp3riA0suWjqbs8vGG9Kne1PrEw2FufVtti58mrWKnaWuEMDssXZlgp+J
QA83Kt50g1V5CzLhWukk4ufxWCwsvkg0XG18sLqAFWC8iwPGgSdWqrl7eo1fiw9zwCz0wwbfFbdP
cBlCqwE61XCx1RonM28EQq5tZoiiHDWt8PiWtgmNH8panSuDqd47v4xr8CT96ey+ccRq7FyBTfF0
61IRx+z0DAxHu0TflnMYiZR063yaTjR4YKPxM2qZsD6QIQaLgQzS67wKKGXTL48JMZBUbStDaOfB
zI+1/LYUjCXW9OGQcplwczpkkX65w9A/20dbDmIeRxAvfycyPGHJ+hxZAKGsawHtZrBK6/08yTwz
KeDklTGeibcLRrgHs96FAfbaiseoTnkd1GHfp4so9IVlg4OtlMSaiIPtXvVLIGU5u+s89MemPNlM
urJm7T2q2/mwBtNCrtS5oo1odzWMW/I3IZA8+9Lb3wu53kYLLWHTmfZU7EpH5y/ObKH+N+/wK6X4
GN3otFW99nzCoUajI/YsjSFIDYIznFtBZu1q0MKy5wj0yqDzHcXfFDsuL+po6pauKsHaUAmFAtwx
gJy70j5Yy4AX2kIpyisVaDRfBzyD4SBTDo1bg92+csImQGGGInDA0o3D5L3QTVn1JHem2X8aeiul
PxmWI3r5WIlIJYIBB2hZLVshWzamp8CDxr1J/rdghurWddFKGhwYArGFsyb5MCINlKsYdPlVPTwl
o3QaE+xc0n2kPUoKzgbUx+KFQ9RpaQsH9Xs6D18/9ZrZIMjLQn4gJfOaZtZc4I6AJutImMr5ZDa+
biePK3v6ZVz65FQzZF28AkQIVqAx7njbebC5FfuuSJ63OB6pipaQJ+pop1igbx38WMDIE+Kr1x4W
9m8CKsqqAc0AvTasqgpRn6fAxoC9fBkEac5sxtr+3Fyga4OaPgVQhfT+xlSl3hV82iXDFaZHmsXc
zQHVoe1TRtXxBtAEy81ALm4SFsRAOOCyU7ZMAouX/USI5wUT/V82UMZzxpEMeSWuLlAhDs0S2SNW
0Fa8bYCRBH7JGBwgFco4IymfUkSG+0wn4H2VoFMc3ov5y22m1cWWpgcRLse8kRNia6jU7H13fyk0
Yzh6iZbsohWj3lQGIYY2rWDo2x1O3Y1Ahdnu/PlzdZrvtVrkx8+deVX1n/y+7BtqYTj+nTh/io+Z
rkeQfgL36MXCnL1wqTJ7m+3eFkt07HXUSSGvxPMBnQ2+JGQwk9ueUwiHfAzbQph1RRTUtguiWGjv
0lxbJA7aHFIPklE0r4pTq5FPM9q9t4mMCP3nS5BHDYQKQR5dK9r6DXHf3/Yq0616oSDgj/USH6m3
NcVzgAxDjEobBvv0HcR3W3Seyr1Li1mFTndoqNQFtpGi7uxuBuoMXqIuT620uNShg+W2sBJLSBMt
fjx2GTbrKlTmrCir975KpcrMRVP2rJztB75e62KULlFHL8muxG0ix7ryWfKEAqYRNob3ealY6x1f
yyTPgOYx5247PviiIR/8ERgR66t2QiKt61D3w2SLYUosOFlyPN8S0whbjH497KI1fCgpHCOsNYBo
3HvG38rkZT+h7DrQcWPggUckUIUK44+RcdWZKp0a8JHKBhafpOBUhsqukl+xaiyxsV7MjfGwNu5E
5MxFnkG9ckaI1vAcaD6wOvWbShtEKcOhqfxKDcK3OVhJv75U0wXjHFnrSkdXAsWigoBLUM05007r
EoP5MMxB2uwUjgMzlSKWttlrpFiVZ7KkwBAphF0APxbbzGLzp8snYDffL4zx9ebRxh5BoylN3izR
ejka15TpVBQDoyV/dn7pPtRIBC/AsTojdg5fuXv9eEftg1nRN4fbRxIzE0pGRTMB+F+o+/aIRpO4
waQWMrGFCA+UseeUOoNu+/iSDpfyMrTiX6CpjupgfiLtYu/kiQQtdEWCFk/HzJUvNBDk7QY47wa+
bWLypzO/t0olMZIACJ2wnG7HU+FbnGLJGZNVnoyVS7DgPA/a5v557su2ohVCoxZhFKUyqslRZbht
1bFEF6EPO2gohRexTrhguGXlO87fwlkWWj543rT0ux1sHlZzRJX32xMBHRsEVv9tKIDzgmyJM3h0
zcJsoe3FraJDkzIE/LnbyJwc72eHB40vPfeFYyxPecK7xNvsiCyS6mecssmOgVtc37+2A2eG4pSD
EmcJQwUZgV6/Raph7fs4Yvej4plEgUxrjubKsu74y1M+6jv+0j05uOnF57Q8s++Chbq03NJ1s+Tm
7cWsBQRb/UuFN6ujgYryS8oV+POMLaIhXyG8Zb2/i48i12Pts5j5CrXEkAODfkA4l7ni8QlOawYg
JXPJN+DwWW6KyvPE/QhxTzxS4978tKyMDe2w6T9HbqLRCjLvxceM958MY0ZcJAA646o8Bk2i+xhL
whEKuw4KvF8hO+llnwy5+w3HSE1lIJBPJHGer6kvw38HG0JHZyf+7iYgsWxBo7KSmlRtSO1XFH/l
i6thBH2lSaSXmJb7qNAV38a20xdByqelsdto5SxqtXBAF3QYvr9XT0JqwddVfbPOHv1F94eoKMEK
jl4p9vbikwR0wPpTVdqt6XIRSeI+/9rucGvUhN1nzfuxehkk+uZf9vA6E04P8uJ8ngfXAGCtM6Pk
Xx9Bz/GYkwe1hcoUMemqNtHaYqhhtecnNBnA0ipZLjsD2Mfwb5mOsJQGATVuAKARyL3OS2mWYdWu
4E1gLZyGZBioJ8ra/oG57XqRLVHDTN3tEhbPWu8VEchXVYqvI61ntiyNsLiHWyksjPkZiCg54+ia
enFFPULagF4HqdN69UBtfShKJ9t63eGgObEHIy4WMQS9D1HHSpNnijY6/NE02UUCRN++v0N6ldxl
VUU9eLd9rrMz8UDbmV5NZajYWbdIwHDohD39XUoeV9+Y1yVJwWapG5TSvnzryCFgNenEaH4SSXSF
preVwOmGEBDTFO5lD06W6thrxaRZddXp3uviFD8kqOhpfmaeWPF5WR5qnaP48bXUUJpv07+dtL3F
GQBnqaRXJIixI/77tlnj+HIYvlX5a1BB4Fwy1OTJur3LF1Bajp5Z94khVbCUKcCtLCwSteo9BuWz
xVF9H3hs1BjM7QLpeaNWRGh1D/6+uuGLhb3BHHY6OnaNhP6yTBd2nYAMhIq28tO1SVLfj05+qwF/
8MHoC3kJh3iU3Gi8eNIdzyS3cu1pH3MGIWxzx9Zr7ePF8HF+oXpHTdj6rF7NLthkvzqhINEVqaAz
4Zzw+gOfRq1qUz0cCMr8DXO3mEkzLDDvbnYfj6P63UAMX+hmffU3SDb2FBXBWZrTNUXkg13Fy9A3
gFN0bZCTCig4vu7ni3QFPOmdwHnyt5FCGXwipCG4oe2axh9QgrA9KXDWTcQqZD/KSnDeoq2WfICb
Sf+rhR/Ht6YQmt3a8LYs6bJl/8VOsf6SVHzB3w3OvXvzCDdGmufwYJT4ScGlIxypEUtDeHxu3DTI
yxArK5YO/pdCo2rKW+dxfj8LhulGOCAp+b/E0gDD03W90kbi+RPNQXSaWOMZRpsBVLnH2ImcPCZm
rs61Xx5/9As8WChMPovqfjB59yNLusO6S8+8ePHTsCjcElqLkDLAwYzsnKlVBR321mv3HyyzT34C
GZMVNEdJcpeV8XeJqXzgvB9ushw0wFozoUzgEf+YUAy+PUHLC9otXMiwcz3QkcJ7Gqec4P5JGhLb
lpF/6QBQ0CxczTp+uxYTKQLOsmR8vi1S34AXKu6P4eOU6HtFRZZUfxY8qTPs6D1qN6GNmrRPEXNk
SXY+u+VslseGSDWcVILvrXdOxpJ57N1VcNAKyMBjy/NUIUo+AELbX8g+YMezZJWIvgQbw4v4wfeb
TH8Bxnw0Ag4NdePkwTnkC5sdx8IxAbuS3wIeHsTOOyx+AF+4C+fdvtJXEmfeb4+CUjYfwewAF66U
fAR7bXU4+09sEJDpmSiyiUBvuJmPjCnIgJWu7TefXHsp+lMzkp0youc3HJM/e/2sBvVtpdGJ8Rgc
c+H9tksUxlgkQ7Wbvx32LEcTb3mbWo1FimFrscbqkGpVfCoLoYQt5i77rgXNc3vxft35c1QMKNZn
6nI+Fq0R83MTwJvSza7MDQzd1V3f4tWgqiNk+1I2kCTklj6LMGkVyqhGLjajoWk+4rbM5bUGgU++
mcA+9RWpfkAq0fJIv60RB6aQ0p/tx5aSv/8gYsnGJY5T01+vJ9KF/Gt048AYtHLRZrv+li7Toqxe
b6M1k0IJ1Uu/2c8E1kl30pM1EHQTYVzqwgrfyjUy6GoMj1XNRNjTxxkgiIs1lUc8gfk9ECoABbOP
YRzmc58E4wjoTpHaosxQTTf8uEDW3G+FiNjnqUvlYW19+Qlit6eJD3NhwU867rLwZlq5ybsmhjEL
cFk3OKJ+3JCg1LzHnhm6TqiULq/eHPV8I2QXpTLadhLTFBRvZo2SObkZNSpM8UV8PVH9UYenB5qI
htFAEi93vttBrFO7vDa49efUMPpC6zpKZSMzqBRBLxQJTXaoFPn/40JRg2Hp67lnMmhv2nQAl1l0
tkQ7xKeDsthrNJop+aPtWijGPro+usg09MOvVb1Gl8pL2aqhtEHPJWE/Hbi4gc4vGtUm4r+25KvA
zstJGhn9r3JNPOyo96C/EbHq4HkeLqtMy8xvmLFvkzXbwjsDzSC4uoss7dez/HONoYCPDndus7t9
rhk3nb9HJxe8wRRmeeds408lVJHV2+zpm63PJoK/rYhrR83juPVGskR/ZxC2QlAntP9aL4WBu42a
sPqdCAi02YiaWove3QfmXqj6jkIMWsczNv8B5SLX6twtsqpbekOyApGqsSDZFTQbq6tH/GWwbJGv
mlXq0LG8UTXQeb+aWyT7dN6X5MtMw6FoEY5jqeOeCuFrSBeuAH6Gzlpy5YKmIvxQS6FhBXj0opQx
hw9SfJD4k63z5k9fWNLkGXbLNswraOUvcAh1Ltg0EALl1GnqSNKETfr9hceNgBj6PZ/0gp2/4Nta
EZ8x+J9SQqcrPO00ESOaZkp498/p2MQAiDL7XNW1uIdMp3tD8aMJbS2V3EAQX/Ia53hditE6/d9H
n/+nhiz1L04AkHIPg/UEhESg0Dodoqe/WcujPzXVLXMuBo/YuHzpgUSub4gVpxJ8enmQYuZ29aXr
RtkvU60dgrKBQjEk4gwaoOMxfR92CA1kWWEOiAtru0CURax7ZPa6Dmd/DG0Mglv1KN+TYjqWNn5h
J89nKFwoYAF2WFJkzN0XBjb4lXpftt1kAfEkR0qy1NqeWiMk2W5n73/40i0af3k6+Hpw7AZlvOSZ
QEzWh6Sb+7MntxUGm2gPxOTaBtNzeHfNzOBLqD6iR3DiS2/+1BEzQH1tjrXlhPS2EHzNBpKbVcX2
3cHrQrQ+CTMJIW9U+ayiBZNlMkFQzUXhP9jr/jFXbw0zHVZwRSx4rPHZewvXUDFn9qv+ehodWueO
8+8Mwcsv8cq0FkIdfabbONTXpEiwBHgsGG6reb0L5jp0StneBjcOO3X6QrsXDtclYk5YYkRiZB98
f9W+MXuPchRjUyoYEE1/pLFyfngg4tCEun+xukgRXAACvM3wIvLi7U/iGABhHa+QmNcKIimMHSvU
7nmBu8ypb0dF4fL21wWZstpuY9yGq2LQZ0wHq7qsEPI7NpVcDOxNMKgqzs3pIcA+ZG4m+377AfbE
Dx/bRhvvNUb5k2kvguV6FRchERmR12vQRpegIWWYvxwFjAHb1nGwMT2qiGLB9pWnzlKLuMjd499R
27SspDieDyMZ2X7xgCiRUyMh+WBuH6IavOmEVSXgHtQhQB11yReAiquapdR3twc3C+Nzz0r6nSyZ
3QJrn+b6tzFAjSO+9v4O/rUX4hQLQTKkWu/FgS2apI6+dx4MC25JaoOgipZbG2bEVIISBSR4aUnF
kPPdKZJkcBaK36CUqNd6wezMezcPIko+FJQLdr8Uh83gsj1C6EtQ9PU9AgqrOHfN+CSHyQEwoedY
B+r8zANWuo9RGjJ7SEfxXl6gwjhjSHxUAfbrU35ZxCyRMMlK/84Jh2MOBGgs+Lb9fRaXK/MgnaZU
xjIR/wbCX3/eopCstdI6PzbKZbpTYrBKRX7rI6vKOb0LkelCSBxUl+JgNAJ/EAIUYrArYE7wQ0Oz
wW8FzX9mkcdR2iQCtVcdeR6Jg3Vw0reaq5ExrKKPvnAj+3veTrr0jJ8UES97Mh5Lsr3y+aY6QbRc
oNphBjXyVoM28ERVFvGi/Odlj6U4IrEkoD0OzIRj9vT5pJ9eq6kf5ybXxTGeDT/f4JHp2XPumzH6
pIagr8aWIu3s5l2nKjMzmTDtX5aC9UXZy4l9gFBT5jXH6h1Xkld4/LlhKKfTH1eJPh5mCNk+zP8t
2Rk+f7VSvDkBpJdxONViSK/zbjuWCPgTa37bScVnZx4pjTyh/H6DvDKUjo8CuzLzJdIitjwm+LBL
VVq57XFXz8CCv1/X9xsikCuxyFpIta7Rcu5iKG2xZld3FhoWTh9KvrTr6a8gYGIyWnmpTIacz90s
+Zy9Eut7AysT/QT6Fh3PmBh1vFyrEMI5YItPRexgSmqpDvYUSk9hmC4+7dND+zYmIOkKM7mmeWaL
69IjbU+lPh6SU+tpFGdpkfwKmxd988rkyNlLz//OlBfqERX+i3dr1svYn8WO3Z1+EDaWFONPcsyM
52y0bFN5GcaY7OZCeVGAfaZCHeGZ2F9OTn61UWMtHizzYxUfw3juF88cjOFTW4s+j3xC238kvtAD
plD7DGuW6NJ+zDVM4qN+DzMIXaTgHMa/8+OVQm7NKu8XQ8F4jX1yrEzxAVjJWuyr2Gi99FSizf1p
kmcDIK+tYEgaNGQatpT69Suw+R2XWACfldOlV8CdWFP3NwWyGCYJ52uZYNvH+y6mG7CyttjAAmVd
kTDiWAFb5TgywBe5CF7vhdO/Y1Vxv8xJdHmSPAt3nJiyAoHd6YtS6RVquNDZGfiJ4V0BIgK9sLpl
hgp1JgflguSghtIup1RoirHx48LHVwYNlJiGODtMKZqAm0w5Q8ySjmzVC4Zg85D1KI4fIAXVqtYB
yIdCwowKXizFE/qcouR6Jgor+BkTLwhwiOZAGBhqDuS4AyLsl5Qe/spxUZTLekk/ZiPh3LXGJDjM
plegI8hZjE/QNjhgBRUQCvHh5Wvxwz8no1oUzuXSYQcjUMDxGyGrQwsW4VvCIQUtBERqgbIZryok
7xQlN9KqUtqTheDhCNtOftGzWlcIE2LRXccMuAUuKcw1EFNhP2d9It3tB77zpM3EHXQvMnHOZnew
uIbCTNRJi43Q8bx5t01OcMO9DFHU+d6Qkc523eE9I7mZZSbvl7H8wpPgOg/2r4RiTfBgcFZUmkiM
GcX5lDr9iRNktMFT5+oedJ89oepfPW8SjeQNuCAzB4qNmubn/JWM3FYM+TmPcyTlWr73fe7OcirH
xQq3AcZSg4LE+oEIgygKgXXaho6TTDbMduNffBeFk/wuF56eKHUnZzH24fM4OlwbDNkxLjFXyTL8
Ce6ZolxyLiqwEn7AkCaTD1/0MrNpRc5W7JMliORlFyAvqciosTbmQw8Ew0Qn8Qlj3VmIdM5F0/0+
8dny1kZ4CrTN/P8RMvdQvQU8swStdiyxDZvHsPJoXolC/0E+XdtSdCDjg/KGpYDp5vLcjLJFA60Z
QHcUWAmJcHcVFvNoBc8CYy/mQYk1+5HZJWgNmZxSYayAlhnwvumhTtcBxIJSJ9LGZdyMJIlpvqLd
Hcx3dYJR0XvEe19yvTcuFwrkG3xVc6rshyMeXwic7H83jVdF12+OTXey02prQWTHuO2cdBP3xTEK
hoAR/NALuBoSjhtcjq/6iYztHJnWylo0m6skLwDhGyR91bsKJh7Sj84otp+fpF/KWaroVHXj8g0g
Ud79/HizWF6grHgfcUD7aKmiCnhDBVjaJE8NCNYFYydFVBFfQgEgoF4OkD8LlIbdkVglFDImDdjA
wpoFEGZWYsfInbE7dvMZC9uge+lmWtkSNczp3VOl2h5B+2gtGl3GAK+xecK24wBsLv/It8reD2qy
LDFAQy2Pi3/ZDHrQISRcPuwF3/ESI/OPaItLt4cA1rZh0z3dwd66hsjoZBT9v2doLT6IpMonqYx7
mmSCfn8MEjbq7RTjVBhN1dT+Izu4yHFhW+07kpeGyl9oaxW+F85+Nhvtgo9yKIr4aWyn7uOiE7nX
celpSGhTR87d9xUDWX7spLFMzy0XAZnM4IoqE5deNzNcYQkRw06hX5Xzw392HTZb8oeT7cc5mIA9
MzgCkqNTHnMeNxqey8GTCyszEBbNW2DSu/clVYt0gJQljtkVRobqw1gHJdCezVRfiLrVnhblTZ5Y
x21e3ueZzYcLTvN0+6AaVLZnfWNsyDnfBYCMxsFAfw3Pwqxqj+SRiXQPmea0eMpl1bn7/eRQBUPc
CwuhcZlV6hGtPlF93RyVyaO4SjyNS6hzNWlbyrdnJ+yQWHi5laywAtXgk2BD3Q5MGNacpSrhc4d5
rmyyvGB2/wChZa6NO+Gs7pTJ3ILBbvXZ50N1Dp3lPiJ2I0pUHPmdwMkls5AeRrER9twI/LD/Z2Sf
Asuz/+kqxkhOn2gBmF5Al9LyFt4P2auDN+weMyD4BVt6qzlW9IgnV/ZFtykCinRhE/IZ0iryBNX7
oD2Eo6FDTtfvaUVey6TEbGmAtRJnFFdhcNguHoIFy1yMzr1NLb2TO2zGKTX/0glgQ6ivrhV/YJ5S
vTxKZKGTH2S2PZtpHSM0U0ShcgVmTZuab408UW1Ykc+/+yQbfCF7DLfB4H47CJu8+DnIc6L/cgIz
0bCWWden19vDqY+qr+RxYoh6Pepm7OLPtFrVCSSxoLcA+fxarSBHqw2yI492+D01nzvjLGWcKDT2
cubieGK/JoAIiiXNZgtd0RClHA2aOYnhiNZehI04vzkwmvXhEjQ4LfXqnHfm+FGpjakpfTMh7lXz
rgqAbL4kGa0Fq0wEWh/PbjIMNbrVgc6PrtWd+ClATWmCW0/EghFTXNPUP2aB8kSmxgsJKrEB8xUB
OUQCMxj42aHB1imGi1A8EiiCzyyaG3g4ZF9BO1KkSbAgQ+A58D1X+iVAWrGzl8HMqkFJfgoEBEzL
CHhJR9wpXdGZvmT5CnTECN2T4Ie+2YMXsKc6BoMQUA59l+VN9/oSI1fMgz9fTprzZjT4+YEQnnDg
ObFra1et5LTCaTp/HXzrOGO9M/9N/Ov9VhvX3OM50QuDVG4V7plLG0sAykfSZdzgYYM+S6qhhdpE
IGxwtTBCttQc8NLeTIBURrhXTkOyJo5qoSDLF4yMxByETWiunUszDstvJX4Y4hWnmZ674FgoZznM
Hkoge/pqRf7JTGGyNgm9GCSsUPTtrT1y3j3NuRfOolZmYyFBXE0x6Awb7q2nQkqBMdSklug4fa7W
jfhMPb7cdkcHDOocX1dKjy/6/3VvrwV7/uzz7LklRm8fk4wMo+2KRVCJRwg9LRgn+U0cSEpHTN9Z
btzWHydOKUxklqWmrtKtGz3MhQqgWF8jKbylzf8mgtAvI6HGPLaQQ4dAnOEMi9ohjFL2CEUCXnOC
oQgQh8f2gCj5ioHF2hkC6qUoq56kBxhxQSDz/pYzucOat0lmR/DvWgW0clZbPwcl2LUZVG1xLgBh
r8xVeAzevKQxFMSGUj5tT4Hx+aGNhFXNlzcu3zDDLiJLwVGXuSGUpANclmL1VDVbMIwjffOZPxDm
jO0WAYwCLWA3Hg6TP8dTmSoKBUBrCVsdOSMdsM3vax/Bw7q3fCOdHzjNBRx/38atqqPjlPT1F++n
dm3c9jDXSmMO6G0jRJ61fXsS6LpvUUMUjn3yo+0+0fjZ263UiXhl4Prn8qM/bMBFjXUbNSEJsKiz
kMlsxKRMo/+vlEfFVgVCMueJLa4svvwcbEiP6+10gZoTW5IjRrYx4pwfyPr/sRov6CnheqqkuT1H
9v8I7Yg8K05Gm2HExn4TQI+18BlaKjrf9fwBg7K6tV/wKcSyleqef3jnHmuHi9tRJ9yYY4YwrMWU
RHt9siVIUiTWea6VW7HgjvfuidTVw/q59n3PjkdZvd9Ji0f4F3k7f7ljvkeTCUqwZQ9SQyoOJxiE
k+M/w2C977ZGr8n1/3NZKo59UZQbcZ10F5DYjDryF2Qh6peHhPzv5n+NoL1A3bKG+7i5Io5Lfn9s
yU7OjpU2FKt3PlzjL6e68Ni/KtPWM6PusG/RCMvPLQE/0VPaxxVcBvXnV/qAa2OB1pSjN/lS3Ihg
4BLrNwCfDctlJUx8KyjqeAw5e9UG550eIraPuI7DqZEuh5VmRrw0fyflWK3EuIP25p+rxMgnJs1b
HlpbM2SoEmIpTnG+wXt0zYtd2c7bBmuem1VzzUayjJtQN7mn/Fv6RbAKsDm93YXeEX3OcsxP3XRa
+nTuKRsIEqJyxTeH6piN8rrQtSLSuYfPir8FFF58Zx6QVPPQPm9beFmuxFkhZ1eBD/X35T5uwe0f
OZJtabMjjanNwEjrJIE+XVFPmzOuvLuTUh4r4rIeaxAY3OqGMrBdnmnA+d8wU3F4JBDggpS6Oxbi
6AGHELT4eTd4yyBmy+xDdHAW2yG18XQtEYNyrLTnpt6XhdxyL19cmaS47ceA7JtzRo31oKexiE0U
FvLyE72DRuW24Zml9jX6s7fqzLYvKTAVzKsJB5taOmNJYm4AoIdyv2aXqrM2JiDF9rjTDtdyNQPZ
4PHOVHGBjqhuWzrbDA7DQlMxOVgDBfOg1f4pAoxqDMF8PlEhbjNIVQzwg4k2+DcCuzMOrsTQfkzA
nEkrFC+2+eM8VmYAg8O+VJxuAOhJq5A31q2m7d/Sl9GwLWofU4J8D19eHKfLHZFZUgfyDpdzaC8P
8UaJAGj3BkiNRARCDlChBB4w7v0KHpfY/W4RNBm8qn9aucusohb/zIaDh1DDfedarA9dvIM52f81
N3BuJmV3O2Gy3v7oyQB88z5e0NSLb2qYP2qiWOQfGlvwlC6fMzwlcH7vEAHj2Q8xLVNzd01CbeQs
qNAKmXjb92qOy2N/bbO0WkAj4lsXEhXHHhu+gzjcH3lqCPt2H9pEXcNr1cASgF898HBWKVLzPN/V
j6OxjMngTHb5V1pSHT1mDxJSowLyPEx0Bqp85H/6HqVF6RlxLljkaPp3x/Yl/1ALwOqufoYwlBML
0Zs64Q8doguIMUWiAnuOCQw3ExFfQ77PgoLEhFTPRpM1B/ghNw3HXdIprgwVzpW1Ut+tUHTGcu1x
M9+76Q7YWyqsa1KSHpA02ZKWidppBxOA3kDMgDYrfjya1hHHmCeMKK6IEPGgJ+5T2QK19beu8Ro2
Pmbzr+DYddsUPWYwMP/A6eWakAp9+7WinDb91VyZeip2yOoVj9FLQ+qrn/o0aF64DKSAYvZFCvG6
J/4Myeq5U1g+Rsa2ISMtRpXiL0R4foSq1zIHo8MpUtK9vR2eAdpIRv00YThzloG/F1L07cRv3g2x
AEEyxd7F8SUrtS7f+DCRyW6liz4jVehmcg1KBVsWjKZZFDbpVISblfgsxjLGLjLnUH1KAg5vEcqc
0r3YQnu7fI78hhaC9CEDCbWIHBS3Dt9kl/qODe+MWNad8Fc+n5unZgbzWlKej7EVL27KeXQAQb3x
4NbaxqxxZWea6EeZ0ojeRDsYVaoM7VBXNX+WXk43HZHRdlEyVXIE9HhwnBxqY34nj368ATrnOWdQ
NRFL62aWpDiESJX6wsn/AQWYQx+lCIsG4JoTG4mkFh5G0UedPLDf59uw5ZdvzZvhyJ7oCdM0ZGvh
7t+MNMzQE6zqcYmD1AjuMSDKYlDMbT3aGEJqQCHKnHU1UMCZL8jH9ZFqdJ+BOgNahoLnooriOYyh
Rpa0sMDoQaPtOqmrG3sp3St1S0DfeCtcaGhmObKJSPu8mtwC6TaPjj0RpwJAn6SO0gp/sQzPoXWh
oC8IcRV9sf9KUNhmO0Uz5h42Z6aremUeRppnTjZ9NwDvE5RYVeIqW370w2HU0aGi6dYSf6XMvVIB
lg2slM+Mz/3gEBTPsYTMMR8FHF1yM8yDkF47njhb0ZU/WsxWXBkZFxi12uJ68DmY7STOo2ZcylmJ
w3hg1rwKAZmNWbF5xuc8WNt/OV2gT7SmCYbxGVL69QuxG0shwPgURHyYywqIgfwL0GrkVmAZVVWE
zGlc+o8xU+FNco8jTRyLDCy6CcnvJ3BN9cGZP6sYJ5fWxsOR4JZUZRWuo7O1JnbRStCebQ+R91Qz
z1UKC9vnuYaIA6yJiXAmDBQbxGNW9lVvj1SqcCxsLcZl8Mrn4iksGCGGTqqTRInGw/Zf/vbIYt1E
URiDOODejM4ipFh6k6hPEWnvGrm81vqz0GTxtkuMyFy6guSJ02NYPkNPXx5JgLiEhmLCuGNDZgt7
HyNddkhr8kPYqiR4eHZkJroCdCnwBapD74MwtWQuq+aXtVB14cXIJL2o8/amvzrD/G0Wms4nmpUe
9X4NIfthtjA4NyRnKSnzICf/XLaOU7wQvyM9wHDAV4YCEQRCkTZWzm3DYSBGuCcAVn579NsoZZ6D
H019ydXfofqTE42v5VWHIc7k7CSz7prlAkGp5OlNMPaiFdrd9j2vmWlSZaUyEkcioQh5AcWj/sZc
gviJg6VTtLUujhyPSt6DKzn/XybRyrusgwMDbICZEq8g44HGpxgcTewGUYMCeNRkdMHsgEd06vNK
XIMo2ZG7nvYyafsHrq8LqTI+qT1iMlnnoQP8SwevBeZ9flNKVjc53M9IXK5OeK5N203Q+tjy63is
rORWaikgSnU5QACBKg5RXv+7ibgAxDiXWBsPJiNb38uUlp6DuSfCJhvOePAlfkTE6yNrGjbzoRP+
lJjxE7ZU3PNOXRm3pUB7Ics2gbTIbOG3oQOYMe6egg6aUKZEUCV9pRFCO0tZP5+FcYxpFTCvzr60
2sOhgIGVtg2rhaA3FXsSJU1CXwA8ZZMObd8q7zOF37AA3LsuJxHxi1u/ggpLP3knYO4X7HT62cD9
4aQZa3kZ5aTG0ocJFIRmGfOowozmBB/Ee/AKs7pDTNBptawmAm++SUAYoZZNM+0wTqxBbm0hMTPt
xP5GXvvE2q+CwV8fiJ9OrFN0YV5fHxNxBCpIQ9IL1DPT3OKAPtJiVaKxL/Ak/51kbxznRI6hDnoY
kmyP7P5xNNlfJqrfenkod5kNBy1I8NyQfHpZTmBnRSoUXziqBlE0ACjuv45O8DVtlJlQKyFd3keH
0HdU5z0S/RJum4PD9zkH1HrMvvYvj9GARcuyz3TdtcP4zFcT6KIO4hpt+iz1dbnHMXpNPqWWoXx5
PU60OGnbVyNMh+8Wcv43IO8hISiY1nM6dpUVSrTZDSxNxHM/J0GOUr34SVp8V8dhxupjt4vzXlYm
o8WKes1H+J2RcZibQ4S4jth83ayD5FmYSX2+Nre8kp293fXssSsYNo1fSPy4j4K3dInQdcGIwnha
W4RJJMlxnLuAHAFR2i0sn0pvR4aG8R/CIyEndnEqKYmFhp1V2zXW0hxNju4dbPO74390vxL8IqSN
nji4FfvytRJ19w5ZK9QZ6mkFm0F8oNyBBqYQnr8gcx75bfKXpJ3+r60a9Dfb/7gaPBmKO2E4V+Y2
RKdZ6o7ImuVUIBysy30DMp/oX7EE2giAP3F26VPV5xC90dHYn72w7UHPmUREKBrvQ5JGyHl9boQs
AIAwnCpdMdRzN91FsgwhQQ6Ec0AZFcUipLp3gGqpO+p3djehcGBEbOQfsJpOtnwj4zuhLU1zBXeB
wZINzvqs3lM5jINkgjUXMQVZKh+szHBfi6cniiQTbNuIlL4KM7JfuSTv1JvfGGH3d7pisW6LpPYt
vWe+HGk4DT/BhehC8Hkp+DmZZIJhDos7scGrFLdpS7L+LLpc43LRurDTU5lFJZ5X4RcSwpaZ8wrn
juvqS+LrKavdfzDsW+cXhzm9PRkpruC+I5osqnAK4lnrZi74gIPavEOcjQdEJtHLD0CIgcQ0INt6
na5rgnfJCxT1ZoZEc+ViZx/k9pTuVWptWSbRTcvPG7JSsEO1AwzJMAzm05yp6Hx3xqDfNssq3JZL
0nOAJnFsVUKmPAzMseDqGWYUAyvwpZxULmLyJiZwsI36TzUQLu/l0MN5EKLaEWrQsIncmLW1sMoY
ZhH3qrcb+Tc4KpcC1kIk6eX1Hon0UidMgQiJvMaFYLRm9NS4HNhzgYSp63J2iajcjqQzli5r+hl4
SbSuEtIHhbw7+ZvZSQ7+TCoPxcvS8tygM84eNGDb6hMN4XcDQGrQV8iWeOzA63HdegHaIRd0rTBO
OxfL9aQEqKExED7qDvT7SRHYls9Q86RZbe5PYTK9TjH9YvK7ifUgiljhFq2d6XuE7Nzj3YfAwZSu
UdYfECCb20eeDXbPBGyZOZbclhjqPT5kl0M/4iThBgnE5cgXzer98rQFh5ecgaSgYj/sV8TUH4iS
OZ21mqV5+HVvyolY/IVw9pBLXn8xaWcZY/pYl/tCHpTd4fVLTpXkd1O4Sn6wgOg4wDBtuV1rxLx2
wCqw+WhHzbbxx5pe2DUolKY8xTRs43dMlJuT2Aqr6LMLRr4TArESfE2BMdvyomHJGModetMaM/Lc
CWEJLYPjWRX5465z1luV13Yg8mDLMcqUMCGBJ/Lx0soJjH8iBXep9QV94HouG+M1CXXeE+keZzpl
T2Nv/ByGoI0hKMj++1Rs/1JGnYlrV2K52mdy+q5/16VrdI5UMm2Va24tDtkLavhyTmZqukWct4LL
oV8af45yZVpKtaNSsyoSkx5wLfMpBaFTjFFlt987c7bRja1IBg4fXQ0DWDy3AHm56RVVpxMkcjPt
Ye0AtUz+w5yQDegC3s8iLJrst9jLTcnw4Ky7BtfDPTcCurPHAANFER1V1OFn2g9Qvdw7nG1Z9QAn
OopufAR3dB/gUAabgoW5FjMNoxLyCPcm4L5DdMt2SotJKSWCo9N93vWkIJnmYJap8aiLpdGess78
nSWnsVyZxSbtPSpXkYIqR1h1aCf0aas7Uu+uj6hHurcB2OduBVuPe56qnUZAke5H0597XkROhOWK
qEp1TLL62VokbkWPzOT2sOoP8ZGGyfgjEOsUDmKDDmcdEoCB3zxHDZNVeVWJ+zEV8oXvqNJKfBE9
HawO92tUBT35X5wVLYgneGn1b3ujokVC+Nizv/l7cwPC9T+3+aJXPrBQpmxIJoElS7ZfGuWiHqay
R6o9QE8gHUrvZAtMgjeNn6xB6tM/ipyRe4PHL02bH+ch4Og4M7gWNEgwGiHNlJlCmQwFTg+XOa86
gjX2WYJNxVuJ6C8JCLLu5ndNOJYcIEWfI58Q8K1MeCAH2TZ5MFq/BxER8mM88c3vskgOK+e4b6iX
ymEEgK3QpTXmNvfx56e27ZWUvzgRhFpdRVzxw4zP+pa009awCQaq+NZi5d2xn1TzdpNsw2Uiblfr
Y2MmrUH3glzBhG5CvLFxp+qXHduGstruGAgJiYQooKxJCyTD6l8ALxKYgBMVpbjt3x/xPkztrAlg
tAjAWcxTUPNLdfUPbBED0oTr7gizmEUXRDxtp4hsAPg2yQeynRMencDURdBtos+x752i+UkjtkYU
i08gRcx8EKEAyB10dGRO1a0oZAPA/Z/cSQODLnF9ALUKGoawRPVnOeoMXwGxQdlB+Y8WF61XP98g
sYyfY+7qj3tdmjU4YH+vyMWCrFG1tQhkteSmLsIkMjYujsDctqUkU62xIJTe7FD66LA2MVqXgWpd
s2clQ3cqI755N7hx4L4/pkr38HNte0niIEzz6anWP4k/Bp6pJSTxSUDYURay1JTBk+qS26J7jgz6
LihW8rH4x4oJXcUhW+hIgSoLlPkLyO9kzWESd0ol+JsorQrOqboxtgodygZgIABxsjAsn96wrA5y
yktiCGhxEN5NJ6QVA6bQrOSj6ON422hBIM0gF88zBKbcZWqozwAyQtjkmupa9h/ESl9rSGBWDkzC
6s+ePSzKUshQ2T3/JXrJz1iY6CUGLiBv7kYnZV2tnIEX523gNVTDE871nhzPgorREDU+kwRuUIEr
vYFmev1j+XJ2B3WsODYzcHzMu+ZcFYr5vP/tv6wvXlF19L7ATYbH07aSf+XDn8jCwSb5mSDewl7l
yraJgoxntkXy0kJg+plOItxmABkCmwH9ZtS0pLuPO76Nn8TkNnMPhsc4h+oIg5P3C9NV/q7W1oCQ
R5nPpB7UiVVXPvQQ+6r5DJh0RzsJ3PnrBbaEA3Q+QLisFA3h5DyF3VqdKVfoEzS/iCbrCdV+o25o
CNsiA6X8tIf5hLwBlLhHZGC1iEF2ikE9OuB+eSVt/D//F4SUFESlnTpl10zCEhGJ+yGDcDYaC2LY
lq7Nfnnxd/iRPJmMeNof4sayj11tZbOqIKafcaRdqMcS7IOqIa7Mx9tze12JK+XG0dh0plRd5ITu
0n8dgIyHtnqet6SX/mgqfWBnSVN0MaG1ODTZe2GhVe9Yh4oMnDLqF0bu2b6a2G0xzLwafSRNE2bd
7yemE7Uddxc0vK6XWfjR2oX/Ktb+t+ERqEBdyOYnWDCl70Lt8e2v0BbKjrIgdvHkdwecNSPzV5cM
Os6FuQIubv0tyP9nsCpECDwerD0ctDUOeSVcD0U8HoFE8Y6TCnK5HtPMAf70gWpOF5PAWZ0u5/vA
PUfxXTskFfxYKxrNZkZj/0a+o8I5np1bBA4J2ZXLoiiD/cdVr0QgSU4lmNFaUuwAI8D/Nmf59/Dt
X6XDZYxwWLZxfnlul4aTKW59lil27qdMKvGjvkTLKE0pcx+do64bxM1amybEYRpRJ+1seQ4KeS0L
HNLeuvop8jVyeHMFRHckcN1Mq8nl16X7uk6G4xQK+0YW5lEYTKbc9VgZQ4tXNFWMqCKxjFMsegDW
jglW+YxIwq3b8wxmwu5KvcPnw+CERn1nh/yYaA8exd2BuW3M/FazPzXU24IGOvqzmUQ+oXjgQX1U
TJ1hvuEM/rxKa6USbKrGxwvb36ajIr87LQNHQErC+cUKh/gL13uJ9Y/ZA+aAeyuqVBa1F9I9YvoJ
PxubhNu4u7yC5sLG4/njLVz1nRclnY/JbVZ7lLqqH0wF40pYx4w9T9vVGNQSZmhW0CtTfk0rrODA
ahLNWBeamPm++gF7SGCR+vZZTxMGQHJQmw7+tChsRaq19gO5UlMUTQW9Zw1lrr5axNQwRJL87XsL
WCmv+d3pE5cbpPdVJ/K/PVr8WkrnTUMHmOVA5QKVFbVBjLGpSx5dINEf1XOgrSGYjTP+Fc25w6Ff
RUbNWj3M1zdirckLXk2pO9TakwgI6OoU1iGEOdzbeWFzg9Xw5o335s4pPDnegohpdDWLA8IsO8aF
pBVLUxY9+FbDOhbhYrZRlPMkpRcOAsm5WoLG+649k8C1jYKrY+5eejzbiWyUf1n07bow7M09uH6v
mX03JlKZMY1HPS9hZWk/RRDS+2edA9w+QLSnbRQomj86cVwUi4P5K2s1luLx4vNwGUUithWkkOA6
ApugzizjEQqR9gyf7LUnBxMoSjZPoRdFrGsQPK/JWpQvaZbmjsx7HrbHfwRjwvXxuVP1U6H1JMgx
YjyYz7ZiiQdoVd7cmootDKQ2pboQ8wwjtgAtg4uaFeKEmyGPqyNycjsr220igS2X1USADKIydtRi
hXqlUG3k196jTxk1jnvLAPqJHInsvl+NZ7FbRSCXcb9E3HMFhgk5aAAszHFT2AmEqMy91mriuMCe
T+Ae4BWY/mvhRpeKdf3vegrruJUi2wMMRxqAJIATrHmqrHnybZd9c9Cy+IWmjMdfVddg5hzFjWXM
arvBzymdGE4BRvDCR1ReFS8LDXTxARjZ21uAxYE6zhO7Jgc3pBp26/vntgqh8HcvqWBG+J0torpW
Rc93cQVuYe4OegIqlacOVTuHiswgUfbmV/TifAFcmtGzNhttt1USHclrp6I6qpkSW0wJimgkhYmB
lrY0zQSAGYRRXxBSgpCwxUaD57su6BZMazO1XQrrnfBl2GacHggFYRigu3bcGTJVAGVmlAPRIVyr
7B3TI9VjDjsPrXj24Z7bVMbGtulVrl09B4XESxPq+2hU+Q9DmmsDTCupwYjjo11mkERs9SMy1Zkk
aEDOAYOVb4+ceFbvtFB/Q7gxdDrxA9psD4ja++k/OBAnDWEJx4guoWP5tecBg6hjKSjLziHYPk1N
WZFOdwVfieEvYK+VJJZoj3DSA/Et2xDZDYBQTt+ufngJn1OqrfFwmGyMkNS7kaShrA4CFLmUZieI
Jx4MckZ/Tz0dSswX+YpoOxaVp7Ex4aQ3624AE5JCvqvhrdxRw5t6wG8ymRwYUbEz4qqxn1r2q/mG
U0pBtkqOUMXFmzdb8S7qgTKzCB5Idw+MdGvF2wapH3YCRbD6Zy++BOQHdF836hXSA4lIYvZzsdL4
KYtJfJTHfQDCBwoU1dc8U8zMHtvov4nYJIC3fU5FnT2tp9fssmhDcwPOliPVs/0wur2YlU9IslRL
e89NZQBClrpdaBuRTn+RAuvW3lIhGr2uVRoGD09mLV9toBIvelEsIpIdj80gi16mG3zKCi4lAMQk
d8R56RdmCLxkuucR7cO34wPp9N1tCwwNM8mKDkiQ/N6yiQRSKgiWLbgPPGX0xjXN90mMMcZyw9h8
DCkfRupB9k9gVzKec+89yShuoqUxpT33GB9zzYUKNVwyA56aIwFI+l/NQjfBcX37zWz+cT5u+iwT
4h5iOlcEiuKNXdQTtnj90Q3iUf1lMeV1+GIKs/C8JgY95BmAZVvMMp5Wlt7FSM2OovH8z1tNpkSx
U5eyP/MSc1BwVi6DLZjgw7JxahyK5TFicG6b62yZCDWepOR0P9N77G3VYZMBw47kzqM+7M9L7Qpx
gJaLm3FDKAvsCBOjhyvQAgTfPHWxI7pa6BoCe/hfk4gYCBoYbSSrwgGcirJlBFUaFtRqwPNpzBux
1lXbgTDOIYCycUloNoWCkBnCBwlvfpxR7CCRkDjRO7CCF3GOpO9skhSwIB50cOPKGISgCKxtylfr
laCEtglVZHMYSY0MVcjZZzDSeeoiVMWEC/Rgog2U6S4YMSomWIp6HHmpXqFt3Xafq85mRoF96ZYZ
7VPjZgPRpgzDEgPsnC4yTExX9lszO1jhrr5m3KQCsSoTDcw6TZ2BXbuLiaroPtY7ae6N3u1jMAk9
sIop7+tshMMk8x15B/CBYZJ+aCkjcZRPLSGQSWbBypEz4HzdjNslP2wsGLKbnrK9PCEEQY6zF01d
Ngq/PhGjIkRzeZtJ2I9B4fAiXjvzC6yWsDcaNCj68xonAkABq9U5TKp5EUThPIZWRbvyLpUY6lKo
GK0YyaD5NkELvw+vbSkgGeSPofSss39ufqG856QBJa/LytjlWQWZeT5ROUCE9vCMMVJ0tlk5bF2+
1dImrPXdXQme3xSg+loz07Fv3N86jgezvOM0ZZ00kWNoMMOsvFU5yQ2kLweAJwSHS/xEgnXU+XlP
Z3k2FgNNYqUCW4ZZ1V3WnRGNIZDV9/ZUP+MJiMRUSzckAyHX5JEoY6yiVsk3T5Ikc7ifhrfdo2Rr
599Cjcb6hRCt0+n7z/upRNRMhv4rOaYSNktJPbkmBcsRH9k5a6rY/4ywW4yRr4iuTVhQsiIQGntz
xJNMfknBV8C9agSTqaY4BYUARK6f/sdPXJGjhDvg98ESGWcP/0sFF38f7WrkDykSPYNeOkoHdxjB
773D/P6vkB22k3dlGBt5XPStSdYPbhDerWWgw0uPZx2ZWybzPpUtb0A7ZXNUO8ovfjtLdfG1M8cG
HGXYO7qeeC3F+G3fWeYF2MuaNj+VT7OGXOLfQeUcu6ner6jS5hH36b9XVMLYn20si5qIBUZorRyb
AZ0pSBwwaReQUh6NmLinIlDpFfwXBVOm0yct2Imu3Yz0ntJO/guzyYOL1zh71FJAwqdhmf/s/oOZ
frkYmqE+AqNNR4OnMilfLQOfqSga7L22OGJlSuoaWoWl2Eu+bC0xwQOgaI7TveIf1OFFtGCxup04
OElMjZqpWNvSOq2vdwpDYaEV8QJCdMu6ZcdxljfwxcazcP6PkzW9NRvUbjjc/znPBjOmRZyzUzNz
xAUHElaY5TwolrN+u5GQW10Hcdv5HuMNRKTrKq2Zg1zSJ3DA7rrkjSwoHH6OLaRpveR4HdrMNi+s
hgBok/clZuQBUuCZXjrdbqaPK6X0hlQosWzO5Vv2hoeIxHM9k7r6glmMEJ2nnuCZaM/uenfg6WmU
IfeRK13uVEP901FYRYshxaWgjYeVLA4QIYp4heBOlMV36VjR0EMufBJOhorfrPLMfAd+MRbhOGVp
R54iVjHi279amOL8uaEhwWLq6ZGdUZcHhIV+W0homhZZ8GGOOVUWGAlRhQ1X1rLnrcNcIwb1+6b5
U3X4J7gAi6UTWI0tdW0ZuhXONcVMcs86sRkwzSky04kA6SZVO5TlW4e9llnmS8N2o818RVmZHAad
6UWmWx6MimfP64cbBVEFx/+TEx/woXGsmn+iaSMhiqEGmWckrP89ijzDYp0eosYPx1ZOXHm2/i5J
s6hl+HOiMiNcsDr0xJsvK3EqAlnHCJvRWqpm+1EjF2l2zi10wnaLpjOrcOg0FaemOMZkfx76aYyp
QBsuoEtJdGQv8p7T/UGlM+IsJ0CuL7Ef/DnNzDFa/1/ar7eaHNLhLoXQ0FTowKLhIErC+4rxDnC/
WBLDrZGw8REYjHab72bdks0GtnK8iL8Tx6WJWLvL2SULDDaOF8A86sAXJINZ0T9NWW/gD6fcQxpa
xS8VlkxXIT++hq95rShPjLp1HLGlxpoaeYAUqu7xvKehdZpNLBPAdTmIpZfHpAs21hNskoPO5xTu
T6KefrVKlLZhFaQn810Y4njdo2p7Lj+t4b87x6MnLS/6qA9GlqLqgF2A7Cv/McVzwFJP3foM4doA
TytUBYCgM2ABEfP/r0JnP1UibbcyRZbovUrL5Z9Lvhf+3G81GvDIVk26RM/fc5rVDrHycGnceZLk
4y074Wbo8XQYG0zF6xuo6mQZn7YPzSn2gh2ychcZN6wcspsOinY0R4ouSyNV9zPHkrsJnVMYOrTy
Nv743lu0H3/CcBonSeA8SYdMRHAmdq2scSgU/uo6XHy22mlGD4l13CM2wuIGSpgHfl4+A5gk3HkG
d3wbRA96aPuyjbfq9k+eKjeHMIPAiVkMfBlIyntAukKHCbtV0OSwHnLHHCvh2G0PPWDOli9VkHpl
EkP6w0aj9LDV27Le9Iek6PL8m/83ScjJFadvvN3NX74t6W6JbFbCDsafO6zTTiz5T/wnW/VhOZ0b
Ja4kh4LtPCc6MUEC/6bek3LNXOFceTH3PyXPRcAO3w25jTId+aIUjceaUXv5y0wqSk0Jz68VUKi1
5XAtzVWzMYUbgvU+Oe8EN5dbqUREiSJ+VtwST1x92+CSv9SIdZNiAYJKTJNKiedE43XDJXCLHIaZ
D+WeslEive27iAl+csXDGfIRo0PkTxuSIU26JwBjsLDeBZrhnuvU6aEWkN3pFnu7BxTMUyZ57Eva
kjy2BSzJSoPevqx7P/1oiUfIj+6MN0lG9v8LNnKje/aXnT9jspXpz7lpFqcfxD1HmiBVUfLb+RFZ
+dIPwMwTG2F2Vx5wIH5aqYPitv74Y0/lXW/u4kR6lUgNK6El3i+45YpevZIVeeb3TGyIInJVTS3U
yt5tCTtZJPR1pRY+tMkYaFmOKlBlr7rGCvt3UQGdZSMEeNlrp7hMdfXWx9pKNk+HgVhpxs6uqAYC
sJWIbMP8YjHcVIFVfHM6UlolTlPawSdHkeHrTo3qwaqIGkUkNgRM4/V+K/ngDOSXeNT6Bm+ZwJsY
IK+eDm4VmW/rAgPbjBrZqhXWzburjs9Z57SeRikU1oWdmuite+PQlXlcETAdsHL8e/XO89Xw/Rab
Z0/b2vs2ziO641BSQnew48QGaGdFMfdGGGjGW7j8JucWmRF6WAp7/sb9nbNpF++EIjjNSUY2zbGF
lKg2IbKAGI3pdsnbTsudUjxTob1n6S+4RNlgxNRby+S8eAOBlDxtyZfQv6YKa594kfWgCVT1G7xB
4SN/UsgXt18HdOuHa5PYqsotTBavHWmVvZCGxRTc6lmJHSKQ/wPkLNqqiUWkC4r5AKdKtKZ+MIbJ
pDJjxdR0BBUD2wDN3Fvf018EiKq9sqZDWX6YcDwidDEN5k2GtJV4vUwuv59d4IV4A7UxlTvZr2P6
cXmG9OgLNM4/C0V+DEAkiOorc2oFo0RjWYSs+SeRM8rDTCXNc40crvwJS+fjg9A1nxdbHyIBct/O
6ikYiFTa5lnFZnMvqePbiczZVAafWQ9JzGZKJVPONHY8PeM5ajaIIAVah3Hmt69DXuwgrJ2SFGlT
b8qT4E2D4mSTbTJaKvUIl/DWJcbE8LnZBKSkWCBsuZ4EzlRpW67orUWlV5XArOe9YllVyL3OD2Gf
Yxuk32fcL1LNgvg0s4P3cr93QPPCgBpBJjgA8bMzp139nz67ZoWV5YeSkAznhnWhXiKzdUZRNzyq
5Pbcox/8/f5Yze2T2P+fKgqCB1VKO81Fr6DZZejE0rmeL961GOEDlGCmD6A+rwXrgO09YZQh7lHx
6MgJSaMvdhURDNJEP3dyEvUL2/AppKe0J2tArEpqVOWdYY8rdPGIFmS5GG/IwBc2sWYK+ia9jlt6
FoZM0qQiHDS3PDQ+kEGDUV99AnVV1Ml1/KZp3Mrccl+sqRXk0OZ0XIJVE6gIfIO1dfil5kT1CSuY
QdGQZONlnNrT3ajrNuMUvxvOcybCADetiyhC9QukYVmmmkrJpOJYYD/vkSCvCBSABQuVGLtJHIpf
JqdGzPb0jWyPvQyqJYqqL6U3wcM0MOgFD0wQ84pGqWCJs/7qyzOJoIYBsDz0UW+VmoeK4++WWm9A
GP8LMHEUzZVC3pVQBZUZ9tKpfhTY8rljpiv1vK2+FxknPPdEVWyYrYmWZXClkjZZDetFdfWbQcb9
wOCYyrRZ1uCNUPkjSXzmjtqpxJa2JBQmm8VoB/oF/d01mJnMuONg6lgRxooLsxjFAfRckr7YD7Px
ISrMzwoU+sblbogxhENS0uXcx+YgtamyTUJwlrUP/y1Iyn7V0+Q5yLLFfmtMWaChY2RWR1psUGqk
CWIdxOCKFl+6PcPpxmP3q8RCoditHNvheS22j9O9nTbcNigvmWo1E34EJZtpn502SnZb+6gXVPRI
2NcOmh+yQW4chO2DV9EjtvQ+Z6Oe9S8uVMXrwbFVDkAN5A3RuXyCGkNT821th4W3lr6L+jAsNMJ0
ll+/rZ2Msp6hMl6zREoYs3a+0AjnQNMQyBXMMtV/5ro+lUQ5rz3RmETvXaGlgDnxxR/kOmZxercO
7j3RGfe7+tSqF8X6dTLEJU55ti9ngOmJk4PueyuN9ixtQimhIbwFkV4YJfgb9I8TGLa0TAY5CHu8
qf32D6KxcmqoUCLeYzogev2PQZLF6X8ikZKlEPS+Ng2cRRpp8pc9s7gdaCmCkHBLlle6ymFMxSUa
8DgunXwr1Y9NuBIZZnhjMIZbZlLBQHum63+g35CDoszgQpVco93F52cboGmgEfMS4kFmZ1M3n5KO
4IHg/0KCnEM55eJHMjplRQWztqxxkXVE4QqXCAMjwZUKs4HyIWcM3VDcfityYQFL8Qw+3om2u+/r
Bk/UrcOxcECP4hOky/T7WfNFt/GSqghiMO5k7oc9UEthBzGriyX/EmGx23/0YYKiedzUqp6pyjAg
TGMx87ZTRG3S92/lysN0Ry2PRzRQ1FjJFzkp4sQdalLpqygvd1eUquwMvF7baRbNnBoXHyx2GTK+
en5nwn6JG4J/p85yU7h8eCoRSFMm/b0Wmzsf1+tI43iZNUzg/lis2GvgG3+RZSxJx0sLbVNT1+Nt
Ktqa+17LIT3VihHVwrOfkf9LDE0J1dsDzTPPzPyXZ29PHPqHNakcZOUCsXn0bxPFM5q0aA03Ii4H
3d2mguIegKGNWjqCUIeFwQs/JegHXDk9qFWC4TEgu1ZTEF3DpvK0XGtugw3izcAAJ7bkK0LHcwCA
T/czc277RwHMFvtdIu72ciOqh+g6zBEfOwo2e6I+svRwa1QV7Qp0baZldUNT5jZDmNMR8dz3iEP/
nvmDKM2coO8EXw70apDLxduAbymTXFsHo7B3n/Dl9auSJxI02Tf+nlKxQNuhO1Z45wVBVg3aR9lR
B0fGYpZMNeECEBRTKgoFhnvRto3kg/GSdfieDmLx7s53braF/nMEZ9NF05YEnNBNOR1YR5WPHRa/
mLgmKVwZQxHxs8yT+uxsf0Exz7L/AVaBXdRzMDjYnZOd6AaWmiJj5FMIAgrC8pLQ+Z21V39w8UdC
tHs84QcUcJgDgBYj75xtj3JbhDZAa8/aOSXnCjeN0MN94ErdP9n59nzg1l4vnXTrVPdfXmpW3rUd
6Q3CLMzrp8TyKqmq2xNjqI3m04juIlZ+1q8TU8eKlCUoHbS0QL4gcwTOtri2SFaMiM/iQXOCxckS
LiXprOnkeuvjJmcl/QbraqKjKLyexhi8fobcTuUzIHoNe0XuFoef6rLlkZKbU32Nduz5ebsnY5TI
3Ip9z7G5DBvhCWwlv9FimjKx9HTHtqXUam+KcUJf+JE+rHH/Sh62r2JfYtMSvIY9UrqXTZG7MCeN
lUcpiGkLSbvoCkO4+9l3MtFSkEvpxh1kIFs8GXpw18580DTFjaPx6t2xAU0HxjN99HMZXgdKGB8l
EiI73MQtOIdrNUfTWBdk1NbNoJMO7uKUtB4SGHTOCvuB8PRG+f6wFYJPiTRj285LbNvDv8p8Vg5/
8aiY84etElDiOE+fIe+1DAUKRmA1es7BiQ5T7OrWF6/TxMG6CKNhKHwLgIYeFWn6NIbYkGPMuKRJ
3yAEkI44bu4AHveOAPykE7KkJjW5869oVBI5AZ6Hu1aNcL0aCKQ2l9Sb1uppSrLCYEQsqJCsMbIS
AkdKxdKxGQPiQ0STj1U5k6qcVg6+OCPqyS0TcKPmVscfthCukjryZJH26vybuk0vgxs4i69LEnsG
yiLXOSe0+rBsLnVprAwgmdspJxVGz0n+1OEh79Iyf5pFAfZLz4rCxpnKeNBgCD9og2GIAcA3tuP/
HTJrvP7LCleUDJKp95wZwlEhRDbYOL4WxJN+W1lVZ+8PQ7Z1rV98JhtYvgfOsqj1rN5Q1K+kPXqk
D902GX0OoyhajNf9HQGITWx8eKioMXCKZ0XpgjgYEMZl2ErCv+jDI7SScM3C8KZP/RFGYyvboSXD
oxErG60VK/wOL2jR4HSD19BTzjlIDhusFDU6sAKNbN2aws5dg/blq9N3lwtlatyIJZhCeGqJlE/O
Om1J/+7hLkvIdUzqUIFXlArurm+Qd6gGKpzlPBJm3GFtEbk0oWcTxUsTU5v5Rr+7Zx/8qhIH9dzw
zXfLbst9o1cZBmd0qA5jJFNHCYIOpxxOCn5LVoIdLmzz4FXxERpWGSxmMMgIvz0NE1wlkPC5pc26
kYFa3EbMH8sXhjwzk15nJ/wzkT8sE1GS/FmxFcs0z6hlIbA5M9skLJwlSo3vGmLOpXFRxvgY9cHK
qCzNVHXJ0LUGqVzJ0i0p//1hl35OyjA9C5eYIlYddl48Sa0lfu4sUOiqCTwvbCgZmMBOr6Yq+Sdc
GJuTbnlF5YTpf4O7ZCeGeSRHAcD+KKsT5szB4k1xkgzuzqJHQZJGhT9BYFT2wkBiOGZ2pWPtF6ow
9WzbqInykBeeW68II2ZhrW3TfBYMu6PR8XAHNYF5DD4p8eio0MTEZN8jsdal7cMxN57WH6LoqK+W
VjkS1pK3KFoqD2YyduiNOAyXDIFXQKqd/irmlk5RJaoTqTSp9qJFWlV2e8EO92xIozPRalKjXR2/
XnMOsNr+hxzpbJ7cs5yBdUBhLPWcOGdhc4n7wlwHmoQ1AwhKNQRyrlK4xfnrprVE9QxcVg9Ydkr7
HPx8gJK+wko8yJn2wctiKCyxXpJJ/NijUSl0vbZW/P5e0wmM0Bqy9NDOuyqHCkuk00b7ULtApRCW
VJ8hqCp+XTzRdDiGY/VyozIEHYMOhnb38MEpMxVBrft+0KQH2Yb6IjZkb/oKr12hj9ddkMqUonQt
92+5RP6rAXt8pMlf44lpHKhghXDsr3THy9H98WRlmcW7xHt4JauWkzmNCu7YqNsfhO9mUzdawsGr
48DdULVNAiQULt8uCtl29Hmb+yQWMVfBYcAwJgrsDbLUGC+pu1LCsQGmrH+UTGTyUehXWZCZOfud
wWcXcTyvKjGrDH8lxQYYAWELzJAxB5VSFAiyE7KYBsgq0lOv6xOEohReG2zajlKMAFpQjCUtkGph
A5D4JK+AIQA+BxmAfCbl0cDp4AHz09IFA+FrSPF0p+rdjp+NqOAa9j1n3YUMg+LoCptxyh3TMsaa
Le+qER3eV8zvQwSc90XluHuhrul9uKPhtECJ88WO+a2KQTDPHoKyjTdlbRhpyZ8nXdksIrXFoi5h
joejUJ2bo9x/7rv+sAUQKynxvFhUUIrQW/RLyWFLEu61J4wUkSA04lG0JBUFq+dUyCh9VgKMZ+Lw
woOMZ0H2oJ+xN9kbhtjMZoSoG4SjaR0Zdd5azFkuRdPyjdJDJwa2qPnEnkJMChxtesaRlav8TgTA
Bjr+ZZbs0/Ngju+JYxUntv6AylkXoUq4c5IsAqnGAD+OHJIOLjb39d5bnnD1Y0BwYH2mjvGH3J4o
tBM7x7eGEPFXHn8RX3Ztb4VLjRnJFIUNmBTi4QSMYTCJ8WUKs1J00fnxIV8Lg8HOcUjAdu5tEnWu
R9ccq68bW9I87sVnba3YeECdhkuWsK343vVN+5ZhHYn5B01ZSYsKIarx/zUTH2pnaASvysh7i1aS
Wgd+3l0VlNR8awPi1fFHeGFw17DyJzT6iZG0WlijY4HN+w5rA8pM2TUWDPKs1zriPrXUats+UAn8
PARrxBo0DnwjxOgLJrU/35yZb0JpvH7sglWHxzMEft0xdenxsNdlS9uO5ZQOSqZD6uvoQDwpc72C
1NPaKhPzmoKyTPGq+TWVehQGJzJEwfvMJN+iX+22DdE8LLpe6G1uKi8BM06EPJxBzFuyBtXEWcDc
7bFnUZEjrHMMjG6pSdJ9mssn9alOgmRtMSKXmrQ+4KHaCqk/X/CUYUUWKvE6gLv8p8ws3QOc0snc
6k5oSQIzaCygDs7067rsEyomNcqm7/souW37QvCrshgnlMZ9s3pJX0rjExF9wCsHRRkwBgFhJMrL
rZDml8IcMbH0q2ymRmDlF177eB7lREg0BFVPWJRBKS0oFClEg/L17iO0B9dX4i4iQ9hmZQNS0e4T
p5eugC1mX79VgFjfaN161x5NJs5pxF/kkvB2vJcJH8N2n23O40gKut1g6xdgrbhot2Mxj3Kox9ZF
uXH45qNMri0lMohOMIf8hmBlKKnyX830lyYnHMowfkiUYq+0B/6RQvgMfHO+0l8XVP2fjfbLXo5h
hseK5EKCIiqWrCt1QnGjtn8zeNrYuL3n3JAvAhBY/30nK/nBpMfENNQGziF4wV+mG8wEP/N0LOAG
tyzep6NmEUm7Nb7FDmXrTDFMCTIcBhyEabZetMwdMOtn+NuC84BDzrNaHWisBADAwIZBlocQH0Sk
7ERArY8YN2gXRA4PuxH0n+dpvcVtI8zawNgUqMqP/ShzkhxnhNTIiCc9pbjLPAmkQbCDv/+kfhls
42vqz8SZ2QJQ/g6+/f2P53h+6GPEJHEhEmOv9WyxPaAnlyY2Iv2S4jcTriTPxT9kgyh01h+RZCim
ouIRHEvr9bjZ+ZduusSX01BnF2ls5LpQytDXy/WiX3Bnk3W+JxtyN7TGqCmLjKcYVVk6Y2+M0sjb
8+Ic0IQdZhVdOGd9QcwPiULMrFT0LdFmZtOdvr/gMS/0RsarjxY/Kf67IkRol1sya/ltaLEbNzvY
2ORKQjI/TqxCBSbZycjO314LjoIHelZdiovUXcgg7YtSnWa/0MqmiDnaeotYiwl4xDHnIyHwrgIz
cgINzvNLcVxGlghc7wIRJKb5j9qNZunv0f1z5MgfKAC+t4/QCrGR0Vt7aoApKL1Fu3OC6qqgUi6T
XL62xiABf5ek10HdByjGoETWaEsIjykEVsPQwHjLcDYxWgArhKyOZEq/YqjxNYCA762xaSMxlQz3
/ZKmWxKfBSWhTVOyBLl6jzGZab1gH8V+5yTvXFKfs68Cbl7AHZLzmpikf31SBFwjkstlowIJUfSj
HLO3yaYp/UOX8q0kUOVuQHIoJJXC6BXkXoKTRgPWECl3pQvFSj9tldMw+sIdED/L0ByV3YaBoae/
THb21XQH9MCZurRQ8dok1OJKpzN7bGzMR5j13eWHgMyk+gC1BhYoFJL/14JcL86bO+06cRgt8M6Z
gSGiglWsGMBQNRLWowhiUtjelploQfpy0R+3TnRta0bhiaMflQDUn6XDs7IAM76nacZngiXBmHKP
5URsebcgsjcV38+HG9a/2igKpWD5vY03P0kiYyEtLkUEVpWRBp1M0Z/WuYJl97vK2LIisR2HgdIG
XMRvaz9JoW8N0tVMhJ2aT+723oqLJY/Bzcs18G+05pY2gN/ngvr8vtGF+K+fEuCeqL0jd8aRRU/t
ZaXMPYuJoDKIiV++rJV/4e2hCyADbY8ZkTAiGpprU9abEyfEioXVe5tvf3DfLUpNNQ7Gho33wz/q
UQAEF9Ymd6LybAujKW3MK0FST2wNLwKWfY2AUrEUMtnmbnSTreDWo+F9YUBR1N09IoOd4zQHbPZ8
4oW4fTqD3J9xygjFtXVYxzP+FsGXvGoHhVDfnIpD4Ow7NnjZYdJd51Ve6fY49IgDjRqINRQBdp6q
+QH0r0mp6uiFBwNAm9JVAeOA5qq+pfNFHUR6rYkqIJzva5eyTYGzc4VNO8gB2RTb/ycazFT0FCKM
rtZAxN6ppSjRPjUJTJF2qXuQIp+GgAyYDgGMMv334JwWuh7rDQqeaU2KUafGrpn80pL2KDkdqmPS
UQSPuO7fhWUvbd2kmblmkNctcg5r/49t+yTlyajb+CGKJ+NUe+rDK+Dipqnyv9Hzx3UPHX+rtIGw
D17XOgENr1J92R2Co9dLRzS7+abYkuF2f2RFPtZQSdC3UulqnNf6U7GmICZT5Je+YwTeVoGI5XbY
imIIfTrBPviqSFBbBK9PUYsUHEEd+8ZEx1AoBysjppaTxL5lChb9MK9otN6/Odl4yc3xCumOd0bE
17HKi6Ns8aeClRs58zhpNrRJaxw97SDBUAtRWsOeSBcxOhMtFWeu3fo1I7+IK0QC8WGWbHKAmMLi
K/zvmdb47svzcm43enJbxlzt7dwf1EggsDni9WTz9F+ouqPC/bQpYyHuKrxEa7oDKN5/uYfJEb2D
qRyBUe+tA4HX6ZwEjUf3zpNdj6gpBxwvdpWpu+f//TEyE+hZd0QMgjOKU8ezQIN2fcXl9c59cpYx
UG2hB7O4JfXdRidz2xeg8ag63LfcrRKObcOOmRLmJBHLNHCl4IC8EZQ7eh5h5prdx1Cw7+nZGqTC
nqRIFLqqJUR4fh57tWs3Ze1VasZ0snkERuA/upinwBLQTx30psvfkqu98Z7N8Z0t0GoCLBt+a4Fi
5QRUgOYt6fdrY+DC8Y+3O/g7udJFlLyST/sk7U0XbXcToBwmTMHVq+JcKHxNRclm1Yf6XnwcHCrX
4w81oQMgwUBR0dqj22Se0WjTGtrC7u94PgpyqED76SCSPE6FsRfpXCuvjZswaU5IP3HyKFnBxHnb
OXSc6m2fDnGL3NgPZh9TEA91Mj3hHh/jJnkQZfaHt7qdGEdNLILzoLOwNTS50BnnxgCVi2O1vLSa
GYK+OFk+HwQEelKR3nv5lK2DJ2YbpovZovloFErfk6DFnfp6VIoWp5BcgxDlSi2XDQ6k2yTZcpkg
po2JVDgK3mhbHx9pVm21rTOUmdvEhMW2wL9dC2je4yvqLlHwnStaFPSD4xVyQyAm1gnQfqzGXJey
EBvvv527MwRyv213McadkD/ygYk5N3T0decL4tz6Mq+dqYH64cIpOUeJAwNvMuhCZXiO44trddE/
D08i9zv1rZvHHZDahGlOFZzGXX+cyaAEPWJw/De2za6t1qEsCSNSZDa7aohEBjJyItdF9PGAYQKW
hfhFLu5bx67bWRiamvEYCrG6pGU3Uzlc1ztEF0S3ftnpThOoY/5fY4RPKglNTW+GIXiSZltOwnIp
WcN6D2LpQ2mJzs/jb3fdtZPME9puJETBDfKvScRyHRp3+qd05m8gpT2lEVJt1xg8K3V+O7Vx3l+4
MTO+LKt5dNajE8WH+tIgHCdhwYDXyAULH14aUhWaWa5z8Ru+9X9TGB7oYp8j3hlL07/XHB9edLZ+
ZYJGpnrIwghP1BB2xZpCcAZ/QSPLQvGJiljyn/46kFGU17jIvMERsv7Sge0RXPKyz01dc8wE41H8
/9fuHqKX7K6eLIz3H3RyX3K2BLcfnMeHlRGiy1CqPXmX5NPtnRQbc6awaqptio8I+g1Vmc1evhj6
xNVDYW+td5vdylcZkjZ3RuJeoo1L4hL98H65OdA4LONBWNqgixxWrcQCcuhZZekhbeKpNT1LYQXV
4pq+fdKyiK6l+ZaClvTsS0yi/SPSShLspfcQj5VcNElpHXCdfEUTXr6SueQSf3Cpf91n0cvwpeLV
ZShj+K6BQ/4OJ9G63Nr2LBCkNNs0eB9j/V5/eIo8WBVCBb+paFbBKQqmHAaSGH5DHslxPpdV0bc+
dntofsrqyQUQWS7zsC2H1QWwpfzzGNHDZ0eKdkwA9ccJibUHh8nqxZPkfspf1O/EyRLGEM/qjAzO
POzy+55Lct2Y9qgKWCmr+HYzH/RItl7qg9fRN8BF3ERjN5skW7fWnxhSzNPK4QrfJcXRqOflnV/6
QuWDHyIYITFvYRf9YrAoIlltQkOSO6976RNjVC+zF/m324daqflJ1Ey97YhPGbssVPC5H8YuJQR6
ne57nQyTRB2ZDKNAsjdjpxlui0l3zadxkw/xKYIyaLlOzor/R0+XtmJp5Nc6qnyXm4C8h79VTR4H
LZ1DtMWBgycblYCm2df3YIevzgPauGp0m3eB5DXsq6CbkB1p03RQxgURYi22SELTd47NuLd0BTI7
8wYahoUa9p6xqiU5miMuPb1MzW4rPU3Z+J2UiW5MDP8/DGVZoA8vOvlfOuNH7tkyyJrh1snUKj+a
RWTWzGO+29oHge2wn+joMrB3zViBH1V3zeqejIdS4ZifeIE8MFlfzdZE2fK2rdqhUW+kKnB/ZCL6
lNdbMYN1H6ww/s9kXYU44MLjYuQr3Iq9GWPnLgjdEno+ID1pMtPSZUsFMqxT1aNh3weeB1gEScAf
zcfT9DwzN9CaGhiceSQem6v8kIKiv1pk9ARvPp5oYSq7qs6TpwJVkrM9TIsQ+hZYrBTgDv30x7Qz
9vcU1egbsMtzeaMH2VlbbOTbZMpQ+d2yy4VZA/c5aMkOYuqUg862jj44sMRrw14pz+cNj/FLU8c2
4POUtepUQwaIH+q7TNqrZs60zLPiIOzMi+vMRtpDgJo9hbP/QY1ehmQ777vIHKNY4bx2CmOqhGPx
CjgpPHRP7JHKq1aZdTALnDJuzNSrbrO5PWNwsvqfZUQE+WXO7BlG6tL6NnG151lnbdc1Sah6lzDS
vfX3d7zRZLnXF/Keb+F1fcztgnLMfMSBuuuIRO9n8IvalsJBKrHXi0E7c5q8MSzCoO7TAY5Kvt3m
ci4HpbTXk6tJ5cd3ixItVCpf/LuHqCYohTygfAigdVrqLDMW0Zw4W2mpJ5wzv3e4cTjvQb61RnP8
R3pJQxcBSpvIZsYorXbZ4+Dx4eH4ZRveNLyLuKZfauJb6mk93CjVVnbV2wn6EFbmmhLTKley1WMD
SQ2KMvFVNy4m6fIL5pwSyZ4VXkFZsecSKDMMBXe0ZxqFv1cHu6etE8gYeVUzDN+rkZ5KOCJpKNW/
LL6UH7JOSa1AdO54E2Km6kmq3yYV6LwgTUl5YDJMdxnHpLtBCNZj4He6AUAU1WNWybsX6IrNS+6c
3TyFFK0MCcTOxPNwHn2XujFj+JTRr7sTXggZUOkPI8zA8ievfBEPLdA982SKGhyYMdVICjWwLi3N
Cg9lCbnQN8O2x2swkkzLx5eaYD5Pw21Muy8SYjyRcHpt8aAsYhpasxkMdOIEQYZy+DDdk/7s3O4/
5seIMiN2Mtgj7el9IWE6qccYNw9yap+uh3p8CDHx0gSzdiArl/390ENhy8WVDYYvb0IDwSHJb1Oo
7Ou5zQunRuNkpf1b7P09JxW8gbi9QFGoPW9tOrqeG0DvnJmuh3RJO8uQ2yovbUBmk+l7UtE5pjG7
QkpQN7lGhnuzqsVYwwnuLCpE2ON7uHYvkl/HvNiMlKhKDFb9MxrceObwDkSTzXWWUSTdsDnf2fn/
ZLDWt7U6uTy/n1z/76ktjYqLj9IJYXa+Pfbo2MGK0VGEoY9C9gutpMgXF2WfjmNaMb6xLHy1xgHe
7Kh7IALlzZ1lW/RxHoCmyFmP9OFY60ekjktNbXIpIkxAIW6j7MGtxx3lwW/yGcsKf3xpcH5kPDJz
mqFPaSoP3wmcqcadlWVzbV6G26PNgfV7hQo+FSxRlm0okTgRo+O6wPpPTZuoUehqMic7sjMrB9ko
0xUoks8a6AKXf+8DF4GMObg+b1ibXf4Kdt9+zMC4eGPm2JYbe4ruQ8B87mHJQFEg+5BYoyGnO3F+
joKhdSgUshl252VWTcO3An/n8JqKUjGDLziepYGC1/1FB9QUScXh4T/wldHlssRj0VUFf6YRCnKL
slBfUEUXprkG+GifMeYvWWstPdeW5SIJa8McygxrGgInrA6tCOzaEJ1prlGMFKQ2qZxLpj8qbPDO
N+vNCi382Kr1lebdfg9pyhwc7wwU7UJo6GEUhVBbGt3IEzwiUa5kIuOfom0ZgmruQxY4GRQb/Ykf
Qk6vx6OuuEq26KijTOqTpy1QKp3NYHzJDsKek/fi6N3+2+gWn9huJGfslb8a9wjDcwTSAv+zUwuk
uJBYxWVTA3BEiexqLFctRkrJdK1WL8x1vPsoDrtbKqf5sPsKkfpPjMlfsjPjoFyqorpYPUqU1Xih
13t2X7u5zhWmtXZlLk5C5gYDfA45qhWOvztGjNFos7kWqjY60dVrKwjUuMzq2PRrfAXXXf0mHOtX
aN8tFrKmfcoV15maB0qeJoSw/SxKXYOmV+CgDJ4DfCdpoJGMBD/iU0/NAgtk0AH2PisgINFayhcD
fmDpF0n+UpAAerkICAcPPeoQ1Rz54OQSNId0q6fFBsth76nOyS2cyijfBCUDmW7zQnYdyDP9+053
wdbiEi40WtX7MW0rWFKPSMdkNLoRUpqJSupxRBVdXJM71wo5F5i31C6T8h31/Lxj5Tvll5BEjNqL
2QgxtOYvKOHEYPZSNQ1x88pDhJzcTNGKDUxU66eBACs1HDPWLYLYp+h7tleRqPls9qGRayx4Wmu2
kq52wBLGTV3q8WdDGB9txDU3noogexM9yW/bLuBrwhZla1SstXd9dPdfWOMb48RiuCeHFTjY0Ncw
GaienGmU/FYQUlgMdS1VoQYDusTYpg31Vj+Z5ZWoECreAbIztk+1oI2BAxJtoD9UEQuneVQgy1zL
WJtWgEOfxfYwukgRSrlGWeRKXSZ4mFmyc4d2Jyo8x/LEIUVAODFl1xx+MQgNZhiM9Hc+OC0fdVuD
68GATe7BXKuWhqvPO0KLq6NbS3ck/B0uuscq0XwHrK9Rn1/sVv7ATFABrXtbENadEdyS5SPjlEQT
8uYbP/CzMgU/gZIH0MCU7CLrSLoiJm4Dnu5//69leT9F8u1YO67zKuiNrOy2buZ4YygPXvYnSm5C
dj3bzM0QnoYpNRPGlPRjYvL0az93NZfGk9g66KpEE+optzTepdoqDIn0cdvAm4ErDVHB1QwPyivH
xDAZsAU9PUFj9GzfHUUHqIb4A75bZzWOkqvSZiWr9ipc4te/rcO8B7+9g2QqvZP6dcGN/zGTf/tO
E7GHHE1XFeRPyGMPuyXJ0wW9L3Nsoz/67cRetbCpiFsYA0M9UmK5/qYVn7Cw0RTMpyOZij4rK/C5
AyZJJ5QagABmuHT5XQsScuQMJrvMhOARSla6XUBn2cO9DSHCM0gu+tTx6nT9dzJNiHxlOFH2gZa0
Ev9WqbAKbNjJTJbRLgZ4zQnKc5MUtFG3KO0EFaCecIMBfL2ON39ZvuxA3PdRtMq6EXfVJxfmaXTj
RXTljtCtguSmmwLhBTXxR8ARD/USFQ8VQy/Uj0OtzOMeKZA4LxCunM++rVylxZkBDVVhyYP5tzdY
BIYJ05rnBY96dj416EjX7HsyZToPsxhMHgLnkLdYsLECti0nfdOzDKHSzN8zHyZTMTL9kn6O86uo
ozGGG/cjjvDwUqeWPSnJcy5M7a7Aadvn8ngpmOTCVBlpZVuXqo+ZyXMoPS604v62BAK/yDulEaP3
zXvznrlZ7IRDEgHrauWGL6plYlpjMp0GJhCk41p+9HjbKFbYFCnfviardKqxyKZxbohP0VuFIM1Y
1e7/CMzaNhDktqetxj/j2ahuQXtEWYF55245Zhv6kvaEBv7snXTAJqU3Dqzxpr0JfEOwBhkEUc5I
EjwoPkPVfcigwEBb+Jv1btsLhZ5Guf1SclYGldI/bZZgGBh5z2HprffyIChn6rtcPKiyp1VHsIOh
QqdgVtT6jhBWTipLo16lysGnsEsXW/2DcqoobxNxyftjBCfnuAtryb1ZFlejAobLeApNZs3nt0FG
qpqfPXmHXHMWnjMt/GdsMcS+1EOC3K6X2v0++ocTAZvSzb4XnhRwDlP0chppNqCppci6+uFOnS3F
Q0ZNC2C9GejzgF+NXq3Duk5NzF97LwRF7yte04X7J56kVjaS06Ty/5d2MXmDoAyriAcCny/ZNhqW
y2Bim2SwIYDp2EPDR9/yQwjbi2qMJazx9owK+DWPCUIUaVE8uNhhl9b9vz8Ygp1UT73YTdLaki7o
2KVP0FydIVhqDZ9fceEC0HAq1550JH2Wd+yuEtNaVQVvFJQ3MXWFc3/YHk896Z+ZEy6LwhrZ5N+v
oMVFEFdZi2P6MwOk/Yo17xPvy7OuuCrqVmnC4HlMPvqWxilLrzN+EWKPEiV0euOcA76LfrzE5mfB
K3kf4pQ4mFMCDD6K5t2VtyW+x21EaAdzcoiD/Xd0VY9qDKCaVQe/YK9Dr/c1F2d88oH/+l2EeC7y
yuctX5EgzVDoxhYRbWX6m/6COeE6PiEeLgiqKiIeG2uLhDiWZ940CWORIX0DFqomybWBz9YxZOy/
J6l7BOdVqFxQO1bIPtdxunDoRN3KauwkWOm7ZgSgUA6mPHs2ipj6xEvq51/L2nOyRHTlA027/0dj
uf3uSnhSK/oOlC+cgBbdErjlVj+QLK+1vAx+2wpfTX6AMFv8bXwfslRgnCj1eKnYQbvxkoEhwKoh
ziT051tDOoaXGhkD3GEWzdWTTgo9OpGFRW9c1++XPxx/idc0VqEVg08bSbMjeb4VkrUtz89V3mlX
jPza9mvoLMP1OXVbYWwsyg+Rm+qTVc6VZtux1cEqoUFmYVwU+ODNZMWnMJecxthbPidpz1lj77p4
ryosewRK6t6Leba7tnSm30UHEVJ8JAvCEgew7Txw0fBsq1h52JRXMA0v4k8+nkRBVxFfhqpwapQE
XRsuarKGUZ+kppBYu2fWqI5dnv7g/Hch3aSp1YiKxlCIrbJofUZJmwyeU2UQhu0wYVERZwwJP+Es
vnoWmsUrQTPOk0tOe36oNs8qWqVCqvEwGnP9UkZbnWnZADzy41fCbsQWL88e7VviEXjuXTPDfh7y
r+VFXfrfI4moRQzw6RSq1xgbftlv6VqoREpeTE7zLwuuyOqY5Ar/TdJC5g0QY0Q8a/kqZ7nPudIz
w7M6bueUftX86OIvbbAEjU+f5/NVD+cnN4Utvy+J6Fu78qu12QYEbBma+SBhnIkVk+E08qYnB3rF
/NaiEQ39HoQAan/FPTqpvaA0+5fqsT/0tFQJATeRXKhZQcJAcl6scZ6Qj5PBQyR0z3e0NOxfsu05
zd+Bcj3iV4NHQVg9WOg9ATQKPYncsw9t+jMFl/FNZuNibI8LilXEbd4vPUCU1J13iCcFJi1iBp4z
a7z3QPaHfouRygGc3nJShuc3gTLUgrMpDHzdQVx2siClr+fMNcxaMSzfDB14iVKeLmvf00YlcOav
QiNzcx1nfFAZ0v7ihJAGN4AySIbW0WoZOY6hGV+SwHsOxDb/Gx2os7zu00PDtM4vwoGoyW1IZsSo
Ns0ihGBw37j6CkhYHqy7fnkWnWOhs3xYn3UbzVVv4uBzDGtfMREFVN4b8LgXNcBN10C1zmjxWkXw
O1gHm7qOQC+6gIHqzB2ZBqTN/WzXS4PgAqW/d+UXjGEsyJwmanAKK8JVOE8ZEDre6cBCB8jmTUAc
ccR6aHeWRuJIXhVxChrqsICsgZtx8fy9m4dBQvGn4/5wTz//ppQlG4qnQhrWJAQFLaFRj1hEOTN/
ZMz6P8LfVZy2N0XI88V+C3njuaSks8rBY4as1cadW8jtv44PzB0l0W7RxSZevaG2fjIuEK/y4GJn
3eJrsEL8HtRrDALKjGumIkCq5qcnOLVOiMdGezMwZFJb904JG9bmomCpfebnsFBhhsf1rom1NWms
xMLGeG95oKb7GxqJqupoP0lJurj0Jgds82f/NN78nnl8IgqwELOYlzYuOi+Qp0pPKzrkET60P+rQ
rDmmItPm7V+1lb6zwLFsXpTN+P9xyNUraULskUv2fB1t0WApD0A40TdCVid63kpeKapw4S7v8+qq
BS95eEun5lzuE3l/ZdwOQTlgi/4A+ItqeI1tfbQUydrAoMo6fz7vtVvBV+vTXIUirwCI+cKQGJfG
QHqaNdDL0xkYJL7qt5FHMZYXade25V+XshrJRp/ifW2SA4Z9XxQy7Ng+ftcgdHTqUFJEqKaUfUFJ
giocjZym1bE79+sHYy8L3fRfFd/AQYReBcEW0CUV8fWEAxPTx3zNo8q9s+N5mMt93oKMvuWACx30
e4bouTrON09YCkFNJ4YhgEw1bBinP3lZyaPgFYFR/TVlcKMuTTYWeU01Ybx7aoRlrm9NqD3wgoWB
WA6z7j0vGQF7lMYebiI1VtYwaV+Oz5L7zAa+ct7EcQzCw9TAfQreZgzkVKQ1KJNxhMEvWvESnvqe
qXwLw5FnbSgYy5sYL4+rsz7gu8Qu6X61+EXrFRVhRfUkRM3YLFkBF2qaRTCWlneGBL6wKuxWeuqj
KUdmSJsuLcsV1jWtOEGBfGXU60llzytEfcfjKrkDFVDc4xu9RLaYDHLIVEZWupPYI6te/KbAKJ49
d6DYbQ2PuPAcTg98w8f8cv4l6CMV5F0GGVwf+VvMRyZ/sZHfAONPIxW4xGfy4bovu+oib37UhUUT
EDo7UUHod+9Ug16h7rakFSi4zhpw/yoXKatNWD63XqHe9Q00sKP4FOZWT4R4o2VMz4H2yvkR7EFS
Q6Zp8U8eane3z+ZaQDKzFjYiU4CoMGwraasyPU6iOYeELtcU9al495MQYrXrm1/Xz4vOh4qXJLL1
X5D0Hob0N1Tpxds3jjzCX6qw/fb3ShxoHcng6I0aabdM2tqsB8EAgiAMFxtGdXx8LNHqMd/dlFqa
cIhZvJxAvJ+yLxqk9j6QSb/NrCjpLjAfqIE7OvWpXHS5wfpc06Kn3PTgxFN2M41eVK3s5GO6r1wK
l89a6Du+MY0tYTec+vMRJc3Suj2sv1GhrqMj2tBN35rKnL+JuWT81FngH4Eqmj5rCVK8GypuLkJq
AGb0ZppEPV/lDb1maJ2uGvAXg0ninSV3tVIG+9BoSBo9ZHNJkP5IrhvILU5vI17CgHIM7QtN6vKJ
cwaFTLAW8pXcIx216ZoqCNPbYpxprzHNpXkDCaJjB8MpWdHN8dp2ycqMT3OAolZyzcTILQ4yRbP4
mK7du/stcJcrZk+6VKZjkSjzkzmJ1TSHUNkrl53idAXJtpWKWLHa9Ha+C98mSvwxPNtVEpP5gocJ
DbjmTfY9R3X62whQv8mWBPefhSS9LpFwt6QqHheqQpMn6v4BTKmhvu9ug+rPgiW4rrsu4L1Ky1yF
DqpJiMwTI3bk9MQQHxIwIbbV76vVT/WCE8WT0YNVqqZPvn9fjiaGykg3DWlgWnco7qBsUJYKJRls
0f84qVo176JeF8wRIsKluIE1MGh9BJt5cXm34r/Lwhv6KIlJLvT5qr7kT8+ez4xttwPnwM0PqTl0
U3Sa55teBaEFt7cnuYRS5m6Zs48u1EaDVke2G6T1mczerAfWZUripWs4WOpsFjm7CPIR5BbSJzvf
Tarfs2i9vsUn5ycRunfOTdAeAlUmd9uQ1rz1cnaWBSlTSAkFlOpu9CtXp+jxXiDXUrPi9G5M2FxD
JbfAnjPT0Yz07KIRv5C4eGOIQmyEMNpDrtxkbS0gH3e+aeic7/jkRW9Zwx+fEcZXby6SBgU9O++d
6OTVXjZhKX1ZRTNRNcDR/mAFPH/Ws0zL/H64whOQtz9YOxwQfZhb4Ziri6ZcCJeOuC7DKoScYo0H
0L7nqZCPsCiaRtEG8AR0p0U/PnCpg5io9UEP3BAO9TrEOvEtw7AaYl9kag8aEPyhZ/5zMhb8AwVp
K+nzhncHnPitZlYITQJPvqm9i/EM46TW45G8KA/Dm4jo93CCIBTMiL9QaQc2e5sR4mavP2miquZU
aiSiCcK0dsyBmScSHS1zn8c3vFefUIvwW0SOKsxj3FAJ7mAZPPSEBIMlUH2ngdP9Eatb5yNcZxGg
TJzRmat/2O+0hyHim/BN0nwuD4ByrBSfy3KZFUuUeM561sPsDlyZBUhJmhBrRb6QLqcXgstzTQ/8
AqRol3fQw+/dOpCpDlZARrzEIzyWY7eXZHLFV/mznvbg6mRd5sHaxMQkcYZdxaFfSdomgYdtGTmF
+yg9yb8qRRZxcxokLzyLeNE6V0918OUVVGdjwGp2+W5ZWhuSvyLuztviCJGqe2QG9+qJxTUr5Fvr
kKD/OVg4yQZefgjaXxZWIIuBNyX6k2VuXt7XKopss4sE94FS5+BrSsrGlYsluwoehQUUArq3nKFL
VlXbf9dx9mMY4GvFF3D0GKhmXuALtsR+bc9l4vlbHocyxsYn2FvVXeO9b1usl4cdUSeGnYkR3lkb
9F9aRcaxxxs8bUa2w81rW3mR549cTOaiVBfiRlpprO0k7bLN3FuHp2mRQMfm0X3gG12fiTpETmEQ
PhqwtfQvePIlwgut8UN23dVGoYvQMNPhwymL6dh5d75puz2wXSvwn6tnRi5H2+CqgXi2UwENn600
TP8c+HOiyjhnZfaDBHHzFW1RG8RYxWWsyHYNLo2X0gxOHUclFTF5EJkVzzHOOjq+4jJVdbDbRqSn
mgUp9asISpIKok2pmkRnfaZ0KvjOoQxoG2F3BV8bOL1kQkPNXTdoPM+ChKsbWqbrauv2p7NqLuWP
lkpz8yb+gO4AaSWOmW4fzlQ1cUO/w6mrKfMIgaaQp9akl1Zp34uDv+wwUM15Whh87gUC6Yy8XN3h
rlO+Th2Gj/99l/m4MEgWWAPoTpeOktj2UlOKyYJpKyvfTiRGyuOxdLboNIHI9l4kK9l+6qQAL8Uw
G04UGlLM536d9f5bzrXZpT/cn+PqZLWwupqvO9kGw+Mk7qriGqldksk2u1R3RrdIZ67/dhSjUHJq
TZ7TiC9JK9Q2lYK8ni2jeBryQOko7D0hbZQZoOW/YcTpLXzQuhAmC50wheuO6r7zgemyT4eujDte
oD0ZNtBaduNsWLzdb4BYxG4IrdDl4BtvSKIB0glQQ8Zj3RDGxYkrIZbOuY5w7/wF0NjApxCZi9cd
CzzOG29zyrl6T4BHA26+XR8vg/UQl7LCo7AQhjyCRXKgtPm0f/2Ozq99FrJ77PwHViYYUNIoFFqt
CfM6tvr3wyzPMOPBtuRNj2lfA8g5+AmTFC1O7pikXX92Qo75Xd457TjcdwXuRjjCS5uABVNKH1id
GRetG+TdDrtgajj6vQkZU/JAUuZpQRTUj1jYKfOcrDZqxc3GlRbIJ+86WAhIJJtEkpNbgjn1b+s4
YrzXVYA5sA6X+kWqMr4dcW666pHdM14juBzMP6lGjFs0078Jpy2azI6Hjq0PpfNxhiIDmtm3z800
76f421E7i0gAs4vgrHhCXT0pzz3c1uRw7BL2doojJh+Mk2Y4qjCwyYeDO3BkRbfWdYrUnPL4nYXE
JnD/NlbHvrrzFn6L9H3XkAHqx1/xUShmkeIDDo7Ny8Py0xkq1fdJd7KNGFJYsN88ASKP9pG/vf7d
798lRTYThBxWkCUfRSzzt1Xl14Pw/3Yg+eO2/MxbcfdNKNrUAofhMfcBAFITqNbLqvjUoBRqpp93
4nS64Qh4wqN8SjqAQRFAHO4mUVe6Y278+QbZbuO1dpwW8U5tYylPdD5o+YVPLABvNJkOJxmFAPGl
tfwYVJNCa1K3K/hGZkmzLBSsBpUUeCS1rwyBBdAVXXgxTPACiI/BdCvnyUooqnVBLwRveqRGNTxl
w9Ok7kJfRumKNMzG86cK3RrT2M1+015D/pIRdkTNURiK8ad7GKf/Ue/9CYrK2JCgB2nZmeeTfd7j
ncRkltVIp1K6/xDctxK6zGfBc3aCfIyb4vjxt13a3CEmksRGvi6gHzcURhySEFdYm0GKGfVu0CfF
ldS7PyJkRmYed3hTxqRpUxkhAzX7kRzmXmb9ig3MAylc8Cu0fkmk47TWJuAvDMCGNlXuf/y/S/EB
zxBIwEDjB5FlZcbvU0IJhWescfROGYV73qNSeO6fECoEnN2omjFGldpVFkp1qdmyt6b++AFsldnL
nFFdd1F2WPxHNMB5fiywaVPSSwArQfSVKJc1YO9jwiufytAGQdPkxlZ29Gddzg0zqPyl9Yw2gVrw
FnFo9+oxlefb1QJp3brl8MBcKIDRiZBTncvI1FU0e+d7MqjFquJ4yd55JlqsKxVS/eW5YQnqWi/7
1n44FTilEN4t53TH1tgCzGZB6NCKBqDm4JSX2DxpEx/FTtyzyHMvJyBkWBRGBOXHSPAJhsTHPfoi
KfATNiAx3G7hO/iYS5gXAGnW+Ljz/C2PPz8I+HKkp7sIcHsXwYIuvmtd5Ku9PbAP4Es5eHtGXLQF
GnzAgf1T0wUCZryZnxXGg8AJpSR5OpEQ9nq+ufkjHhHV6Ccz6zkKsydYkJogUeLVxA32wGof4pK8
kJ5FRK5LV8dHD95H86VYehAg91X8klrVBdSX5dN+Ji7L4sMSAOckZbkquWUDgonhl6zXB0LcIMCa
w37wuu4Y9aY58vqy0lvvJg+ZJDdt+525OoE26gA9N7t8y4OU8zj50cheQwabqS2x9Rcg6T3GBzYA
DLKhGQogPb8dkJsdAPP/jTn94lCXsaAXfJtSVkfrTqpuz7CuWxO8hRUcIQqhQQNymeyOx5itMoND
ruzna/SNLIsH0suL3BqDolKUBXN+el6JmKLIjub1oun6k4/NnDx56NvbxgOlr5hR4bPXa7AffLbV
7nNEbDC/25rcHVtB3iwx5VMZrf0Tjv0RN1spAruSKkae1OGFYpE/mR6VokjjuLsIdoWaO3BCQloC
6cncQp7Vs/oYEfMUS96XNsWbOWXokGKvqhj2wVghntaqgciQxbRGhUiW9gHNkcowNVdNOZ10J2oJ
IufSqECvQxGoTe+AvaOlcd0xM16yggMKA1WDB0WO2qjOUzQSxUm4TlL/3tz7QR5oBiZfBq1M5QDT
vIqs1WfWb2xoUF7dUAun0/SudcTWdiJmIvXQ+udv/eMUtY9zXo3u8j7ZcnYzFLq9tNpVa8gVbRiO
UhkMCQdald46OqDPhjxJHqUeGNV9619dA3zTY1cP30KWgtPFNT0wtbup6s+NRQJkNgdiTw7zbBCN
o3pabW5mxeWPb6m7EiKUB/Yy60yBbY7c2aghuWoWp2A4Oo4SFuElELomidk137Mh5Vun0RAminq/
6ExowdmdcY9oOztfXlQEwuqRJQKChnTqKyfU8nN5xXTa468ToBDxK8iuiIqAiEhYPW8qEpShwdg5
EIT1HAkrvQBFYD+wfMOq5C8ZExxx+oXce5bCQM2d5Dv7Vsx2qjL8cbWIeDD0DNzZuqGEgjkYD7N7
cV1z9kOLOLW8+sJzXLjJlQKn+3ZXQQ4PVVEF4y1OZ8iSED+9iTAg1ynIyVz0Kw4OXuck5uHTQ1sR
6ydcIi4EeWLIx0Bl+VFOYQUierDYkDr6HRWeTOkJidRFGyova8XxjXK2myv0P6Es1Z70qfFVDIuU
yA1QL1fdqdUIiYHIQLNAzGeKbaYWwsi4DWn80I2/Nj/40BEVz8ZDDUmBLZ59mw1HSSgLbHewRfy3
qbEETdtQzbMiAt6IZ899rzFmBK4f1nbi21YLfqPOdF4443DLOqSssu5Mw7ZCSEGpL4thbBsDx13S
+AXOjDb2ciL1GGf6aYwfk3NxWAIXO/8XR35MXcQQk2Z8v1dz3nQvGx9hrGS5Ij37uY4IAhVv24sM
BFK35ZjRoENfvs7sNuq/ymZezC8cgk/yXbzNbrqMvaeYzH/44WrMosxLF09NGAGoyUOjP4TGHFJT
89DK5Y43El18tce9csnVTZps9w0lMpmSRUsCxsVm7ITBS3MuZRRTMmPNNe+I1b4qu8g9mXzMYg3A
rkzsUOSPdiu4keDiz0vx5P/tEXpEIpZp0N8qXwVj1gjvUj76454mehDu4T+H6iIz+OFhIU4iFW81
UjXMTWkkZtZk47YMygOJ90DwlArR6ipO7KYnhGN55Pud8YkPg4/ow8nTKGmxiUXI7YsetVQfLPWR
hkQ62CvlxPhy4tseTQdmrzMUPomCjcOlGJDuMh2OwoDfDwalAD8pmVGrCCKDvduJHGMopSUDIYTy
VCblzzdV7srfATRIHvXY57UWIjqCUAzRG9st1NoZkxhX710E9iOpM0dbkIYwHDslacVC3bkcnFwY
SJ5pAVUVVNTWr5R2MYZgXkscKOV0LhspKVN/W38HP1ZOVCMyVZ3UyAs5l07zou4jYEGgWQvkJzz7
6qJLm9+2hmuQRCgeGErv7p4oBi0xmnJXjGW1ToathcMSlFSqf4r5dbfxRrACt2O4EfSoUD8WmHfB
7xUpcRnbVIG9jOOKZ9bktUeeA48he7l1LTl33N8rxQbSKPXKG+TJpeBz5P2FEuMjS4DgvK56zaUf
mPq2bExovhe7I0bBbbUCtBR9F3L9slicKQE9Wtm/Afu3q9O3PjojtcE/Ho7Pch7P76Xuy6xvFXLj
6tBvf/p5ZLTbdnB9Rlo/ngo9wt6ot0xzMpEoLn2lbdAKJu1tpdQ429Mjr1mZedQ/BHefmTeKWIJH
CSufrovccyh0Qn1YSRrKH0Wfq/qVREn1ULS09r39diO7/Z8FwOLK2I0RmEjnIddGsJ8fQVpWe+iq
s/a45GWMhi1qOqilajuDxIu8lvPMuMTNHmNTg93ALJ/yips56AL5aSS3V2UieL4NKZTO8/8JwU/D
dfN/k0VULmrD7LOSYcGTqS7Yhh3Z6uV0GMMayHYYdnLA3943+ma7AE2nq2QLm2L/gcVBtvhSa0aa
F6jP3k1AcC6GVwfyVVmk/QPNzkU7WS+vrI05GVY2k45f0iju8+l40uhlG7zjjpz9BBMqVmUfsq3F
NbBYss8dmX0dbj1nccBa4Cw2L7YahbFx0kodBxQaVl/TrE+TccRDRiO0BFNfutwV43nAHmROJ2yL
7iurZpomJAqMMVBYDDCq/QOeSdmlYQP3/0Ex4SJOFyZtEIjJ1+X1wYPDkzqGqeLAalOiG7z9yzPa
DqxuG2cEfQTlMtg9GAN9ANgOr/xWfhpmQf3qUzG61rkildtdpoZQUK79MAUD6pxaCv10lagbBX0O
dfcf5wLjiOGB3Z0T11pzAS7SBeRxCAsXn+v2nmvEOFZCw1cj0BuUOv2toS+mJpEjk0gcjWwfZpAA
A65GIMTg1BqdGqruGRVOsx7ckSoPFvTbStRkiHUvpwqy9oBe3r4tF9t6F7NvieOyV27rR1Ukg29d
ybnEy+HBe1Nse4vEvjk1B4Qk8DRYk3bQF8G7eWgw5k2XlgzijNLh2TGQORgzem6/AyOwwJaUINuJ
9NlxbDupDXn2/bBDWMcUu98mDzMNsLq3gcsuCAZwQ9wd1A/e7j5FQIDl6oxEd2H20ni0f+B4b7TC
8CUt56lwrclPsvemMhoEyRqr2DoIrZaDdi8JJqESOcY+wmvSMUibfrXnGN/HImqI0xYPt2b28qjj
mV7iYB2UNG1RPDF7JxN9pHFTYflivgkwNrsWST5CwnNw7Y6JO28sNrd7DeEbzQ6wDhR35K4Q3Bmo
sBuq1T49rPpyOpAsIAaEAiCY+iA1x7WLLY/QMP5uoOBrPHdfBUZm9MkNQk0i09wfG5t7AChWlst/
iZB7bLztAlqSQdbuwc6JHJX7BQ1E2NMOspAWMBNHytHfw7WS3JxBm/+CCsaihndiQo8UJL/Cd3Jf
Ilz+JyT/u3lgU6z8Ps+JokyHQSozz+Chtae4H3rJ9qfeLS7fBifISNFn363L5WE878fp/Mkw+22n
wj5if6l1QtslZ08l6oH7AjcsnP3s4S4Rh0yTsHJZaWWNJ9noJoqse76LwmOFBu9RgwIfORm/rQjP
FqJknZI/5Uao7WL9ObUnVWckJjnN0RKZw9tbGFSMIbjFkkAOMdg43LFN87A9lTAMwjXNr0kFTleu
FhulUQLU0qx8jwxKZ0ixVrRl/aVoYC29Mgt1kYtwh55FbLEde3la4hNFDE+WjEHhpE+OWdX8qFV7
rfJYgSELjPKMMsS+vzzr1V6nyTIi9L5IqRZN1m0DJYT4Di4MNAh2zLYhrZozvIkm7pRlQisTQmFh
4ym1lLPMMklkDIV7CkMhSMGx/VsqjDXpJonlcXYwKGJd64IhHEbwLgeyGbSBdx/+wX4dSVIldV4r
K7NosPcutu6PEPI5tXPlFuXjcLUA42JjbwmtB4WpU32PxY4BOlVPOOXHvDnKJhNayB70IC1Xo8eZ
fVwFrj8EaMUrBLLiVl6UgNsnggkL//DCVKXsiiQWefLSHFug9F0SF74w7n5EgIrRAtmJbG/tP9i8
pi9GYd9ImIn49RNn2rGAg8bA/IPagNwIdDqzVGphPx0AsKse2MtXla+tlPAOr1iRsMQolvCHaObw
B8//IJPzEZC3dASQIT9tJIvt1ILV7dtjjP9nU6Y/Me1KNF2kcUImwvupaSy7nsf9FOvBy89yJHNo
lLjoo52VFNBbdz/l5hnMwugsl+q4zsnrlszxmYaw+vAQbgW0c49VZSj2ByKvePoT8/yiN3qNoFTA
TM4ZqEtonMD6ww/ooh4g7DCfaZ5KltgusK9VVehAidbml62yiSTW5cm1TANGgxOtYTCcKajOQbk2
+gzYqIzc42hYETKp6Za8jo6EhZtsdNPzzHyf5ZKDFVPexDk9yhIKVSVNcXW8S3p9NOM1iYoekPS4
VypQImUk94rp7dlUrj+9FfR73wsfrxOcx1ycietKBxP6RDaSh05K2rajETiZOu7MefcU7P6aV13w
ieOca2TyJOwFMskKFoZO8pq8REKiGXZ/v1d/Pn0cgrE6UxB4hmRFKhku2UJxyPGCcXH00bdkOu32
Q4jjt8E2JOxeti0Ht64vtBTGeUtbgNc0HEPjqS2l30x/J1Bds96pJrtxdnHy48tz6HYDXGW1Gkqm
f2jNpIGmukvNwDBuYbBH0Yco77hxX799uJFJFSIRDVvxUgVZuzLIN+LvqJxHLbse+QgaWQ6YmcAl
STPuW+rONN8owF7B1LwVH26GhP+sGO+qZ52dEvUHrZQMFtxthbvmepRvqAbqIEmhnT4eX5kWQdqc
iZL1gpnvRbBijfj1Vx333VLHSz3+B21NYEYC2we652AulgBbmmUDNXh6iFcLqYYwt6qyD7qdpqDZ
urqnwQPw7wrMvqMShHvxuhY78IminVpB9g/5JC3Zla3Rzg9XYx8Jj3h3B9Myep6Y67PO4bZvpx2E
Ejm1nPdMxaBGQmuXjlKSTj07/ak0BaIGVayN+xB0+RtLNnZ5NZEwaGpXPrj1GlMqBePgKUt+pyd1
wQVND507CH9Fv+0ML1tU0Mtbo+NszMQ8SZWaAAy/DfDkO/kI7qSudXI5PLfGWvyGpWq5epY4A7qg
pW6ZEm+5rSyvUP+ictce22BD1zkECXrB/QaB3IwAMdgmdV714y4OozGJd0DNVHWk2K/Ls8ev5JcG
XpK+rIIXxiWTCPl6S40ysvyfgFYGb8sKR7pfThl4zHegnXfzTj/wAOvq/AGOxM8WcBXkfiEb9zGC
biidIr0LJ4R3aQSZp0EWIDd+TxI3F+KwOjvSN63aQhvaRSZOFHWwnx9RwS93lGCkqVPXHpi32moA
vWxdCS0ZbFp9+e96+Br2BDleL1yXvsRfKpG72BBBHaYWXXvs7ths4tu3Me7V0H2iU7tcdOBMnvsF
nkI2GGHYWDyH6Bi5tOomj0CeGBfkCQwhfNcIJ0epSFfT5pjQcA5ZAdRvf8zCp/sx8a3JCPfC70+W
IvQkXzrQMrBLs2oVBOsQstfhMcYC/JMrtl4f0fN1Xvs+qa/iSekRKn2VHAnltc/XAZ4/YXNzushE
8gJS0ykNXdzAgPgVjuxuKrD5h5JNuo/pPcr683UMlXTyZUbaB+EUKq1DSC+76Uh5jIuDsxisySsL
vtp1XTbaugPtp45euab5TaRFDqNd1kRS2oBiY/HBJtjWlcxvflKkSIKAPvYUF9FW4GaQVVVfjwAP
Fa+ervp+PnCf4+tg1SFwpbIOpRIWJsR19gxM+FHRHS7AHe/lmO4pHwRC8pKP7y5fpPKZPofeu1jj
rbWod9fYM3raAUj1MXby3C4ULVgM6WmrhpHzBZUNUvdXXrhCsuKW0I9isgahcv5pHoNhHP9cJQZe
B3IkqUIfqlVTjN56PEir0z2G7ntgJQbHtIAF90lu+ZM8WpJ4brX4sJwvpATU41cV+GVedsJB8Ajj
DvKXbXO4xQXR7bv1x24jSCm0TupKcm2SQmIWy/7NoIAxpVeb9tEjPF6/J4/JJrLGl9V6joTBKT/J
Hr85KNubPWK9DZkAOEboPwxNrqAQjKI82GREY5QLeMqTUc9xxU3+r8ROPydzkPObxbW3BjmplNn+
K5oOpvieO6uKfPD8QLWRHDNQgLo2ZHGg+ul2dS9ia9WzQjJ7p+Eh+3EH4M7IFwKYNI9XxKq9RRdu
ATXng6JcWTXPzPu7EJ0aorcyspfvUAWdVcjHQrKcHlB95IJvWlgDZQollznlr7N4MOm+dO3Xi5uH
i7DX+zNP7AArW0J2IfyJ4bZsKPetxMJESgwSOXmyZnZ0HmZq0jeKof0em3SC0X1xrCuuFGx9WFLq
P0kuvq0UXnY1kb73yRI6L+WUgelxhGNCbseTSQb9fVg93NFQdORcxF7+D0a/UM+SO8/awhDcuafY
Z9sXkMigbE3t3uzdbgCBBAEwSMthi+sUvM9r/SG/JGAfko9ezD4x1twqywjfGyOpYXVsXI6D9U3n
3BXcru0D/3qxVlIbo7PXiI955C2epTLE3Fqoh1052fLwlMyFxEBAESX1pGzaZ508MOxb0ylpESY7
L1FtDwR5yUt5I3IAcLKS6Ge6AHlnU7iFdE9wjqiEi9WD0jpjOISkxnw2X4z9gnwFXi6hCOHaTl1L
WrVBvF91iVkSWC5Nrs6Pab5E4EoZ9JPtmqQ13al5M7P+u9xR01vkcflCN2w4J8HrYFj0QvYFX3xR
56C17IcLh8+9sI2ccPwWKkXvKYqvWhiDFuB5+iE4ScMkQaRp6JQnaDIgmyUZp5qE/kqelF1Gqyts
ZPeBqKTiYVkoxF6msue+kdJZYNz69OBqb/7uYmUEHHeDAqRp854D4XrXsdAe/j32D13uWBdEFUxQ
UIlkFChru4SbR8IxrsTngCzrO+19frhpLQqT/EJ1/wlCejDdG0AXGeDn3di13PTs+AB7yEClpgj0
WYVVItQcTpL/u9fcN2nMnJqpCSjkcDp1Ks6164IJE/HHYpuxo4OgK+tV9K8AKPG6kwm03KQq0BMv
1cGhT68DheCjuf0r2GEKyOzQYEmBdV40MC/WDBLL5hMYMwiXxeahUj8DWRE8jqMV0UWZw9gJt/SJ
zwUcA2jDj3EPsybUezuJm5EW3DJRl3y1FWDZoSpvQXpcjLIEZN4klmLt9BQay7RspOycFpSGemua
OktJu6hZGK0ZZzy7cpCUEFhA1naKffWnfow6kXd7NgXDLffzkCwOjEtgVVcs5QcqqzV8aIibvuOu
YQRxqlS6oxl/Bjn1DQKdEwt5/BD5dLtDgQSCFODptsFS7npze+mwlM4tTPy+/lO77KmjXK4WdayF
wRn/wfYQP1E1nZrieYjYCgxztjC039xWvRHWzXrxkyW5G3ybFPks0hb8C2aF6Av4f7iEeWOpYB/y
9xWUMVz7ApRmcKvdMH4LgAMbnyh5jyMf4V/8F6MAX6Oz3nU6Jd6weQ1etOPvOxZa+WA+26KiWbVH
qoAcPFS5V+uKPbQag4GmHbDWodeUhjc/tIFMdsOTvSfopdfV3xVYTRNJvh3UonnvTAtulVqu0//M
LYgZUMH9ddOGZJBGyfI7o7MbLOABRg7AL6y0aeIH0HwTZNIJgQffv22gLZfhaY76bu3j/JhJjEJZ
frJhyELlCvDHIsqdTn+qX8FfAV6j7eCDGhrCr1Y1bUo9lDIp9eDQJZsfe/ue8l2iWBLspp9836I6
rCWzkdhyvVftr75ttxuyMzGEdVam34ottstp3+trE3c0H2wFH8sUbQj1ZYFZiOYjSZqGpXN9EeS+
qjNVHA0V83utvyRAtalXYipeXps0xt0wTv6dTHwWnv/ABBEGVWa+Qlqj3ruVVQRQQeNq+4N9B+sw
V+Sjvjn368NGfmQfN5H2mPBn7S/9egoMEBLG4xEcQ9Iv6mhyvnx8AskjWOixb3YC+vRLWY7TEYnm
8OL5D0kYh7C1onYW7XfyYQni3xZ3B/pXDvHV4zo1DNzdu8YDB7gt3OSm3vXwW3dJ9DWtxNFrmSS/
4fcgwzc32KdU/qO2+iUeAX4OkxrehPpzzXdeoYvbVtE4/9u4O6Qjz4BWO/mXhPK0BmYL3e89ALxX
Eib7KlLKdmzCr3TyZ3fPAknVLYY5GpTiej/qi6y3Y5qgla9Fq75rDO546VexPH21rqKxM2Z6USgB
4JoikM5xe4zCkk3LMUxfd6Ei+IxJYG5PIkym2fN/ybvGdNK5D9vhRyR3Mmwny8x0nACa1lRAdKuA
Y3wswFYBA2Ibf94vZaxH8hhWfLSVvYKNQJ5uN+nAIPdlHIT1+5tAJMW3KW/Eq0t1UX5hlutcA7v2
adL9B7lF9MFhz/8OtKppB1fSCHyRacUo6gLFf+ivw0QvMUk+4UAtDU5U4hVcCxchMlTledkFRMQI
C5MVM7803urfmLlkLVGH+jkzUTr8iuqBv+cWUZ+EYYv6QdA/uxintxrtKGbTEMF440j0jyv4vH1y
vmd+2Ji6pQJRmGcr8n9d8pvupFvNikcAuXM4U5uFo/1H1zg7qQxWuDEgg04FvM68G2V6DPP5DPah
GXYUlYeppGqm9Wvi/gJ57WralU9H8CCbqBdjJGAbCZH7sC4EQHZObaNftcZr9pDv4Kyi7kSTIszU
y18K8AZ3+5rJdu1hHk7GFwVtB2FtDM0JHvHKzjvnL812ilOnfed5/XE4MKE2i8dL8wb8mLVBDoFy
uJ6VIIq4G0DBkTno1HbAbRF1GNIbTh6AWa5fewfEwAtv8Qo8AzSIZvYmvbYeOAq9afJIB20F4T7W
7JlhhiYNyuAhQcGKCsN0a4oKw8QVHHOKm0Ol5bQBdLJsA1AV/C+FMR9GUrgQ0CY2uWJikQqZpToM
F1yAsqQx4VbaI7pBvRRRLFx9E/xj59nVCROwJj5aZI7u8ls2LJ329bQDAcwRMRv/eH+mnU15fi/T
MzA/NQxpd2W12HXvr8vQCvJDCrekFmuoJWvYDqfOQJFwbv9gEnP132IxrkjNKbN73qt18uYy8G2V
2I15K5vlrjh4rOHf5J7X6yz7430Rp407nDtMBCZHiPARO9UYmIeOwDbFusG7QlfxGsEekV/26fM1
Vq92L+1HFr/PCJDPy+3EQc5hlUrRU5tfdfxaXnS4qOWvPmklBhrlbNz/2ZGp+Ao0M4883Gljn57v
qIzNwPx8fQudNAucFCXRfTw7x5NgUne/uJ/Jpt6lrKruNh5FTCvwQbKbpLn5QgHMSYaJFC+qhYlo
YN66T8HujKgmcKIVrebyB78HOEnvXeZgkB8nOVlUaqeavHh5fvX7uAXl8/nDAl7/WSxy+mNGIS16
CEiDvQJH+JcecTjshhMTOX4oJYg0jfgusrOrURuEwLssHlSSqwNXvEC3Es/+fBLkk1ycmBAEPsCa
lD7+TITEiyJBkemNAdAj9rC0tP7++cAeuaOqSXS48K0U1KfT8rCA3v6wTvHRxMqnZeu4rc06zKiE
jauyzlQ+cM6DNmmVn86fq6YZTge9xnMr0QJdNBRixmS9nrZE6dNz+VO1BtlhmmaL3LiKiijLeHxJ
wEBaCCFRKcZjALcbijjTnTz7C8Dv0P5dW6Zx80xmEmTlzMudfjTcZYHWv4Ughy3QPh8w1W7o6JRN
PEB28wNyMjmJY4T0K1STmDdGfzCLZpdW2yQnmgQakntO1HdysA2Vt41QZwKnnH+wR0FYU9k60CpJ
3ymYVJHzO3dpfTX0mTr+ad0U2NDebw+mWOD8bqigsc70Nuz0bv2hR73+QKKtv+wv05xGqgTV0Jnx
1HRMUcIl3poKo2oYRMcglzqV9Lsng+7DoJCHsko/KMfNkOVnsAfsdcRhoyU/UHpLJHs841G1dyrf
WGDcsMmwJbsuSivaRVCBHv/rpdPZUbOwtaNypO/elmVHaNF9ToOtwJ4r/FZxJhhCu5OeXoKk37X/
nCl9TcvagrR8XzSg1x7UJTnexDzOErrgeX3F3fsWWllMlatoOBMdppbCbzh87AiyOIWiXrrRBprX
FqpnzzBIGnMq8CrdD199EiE787xQr9Ak0jnB3oXl8pp0dja42S5iZ6SptQvrlQuXDfgGnszLxtrB
WwmSCM7FgoDC2XfpDHtVfSgXhltFT19Wtwap+lk8EOQY5HLa2v6MAguOANTaAh5onR29ZMbtijxH
/HUGMoHqXFxAUofRnF008XtYQ21MyMQKkdWeHfaXFkRkvyjAvGqIXUY4yvn0qJiTm8pqu5hHLsE7
AmSsl15zMHFzdZQMKANVCGPCOFqU51R1ilV6mqN76D8HbsaImd/c/TStGYlhoJys6WJzCgv7BPLF
MOGm5ezDqA2AnfCYuYww9ORCaERpBmuTjVwEwTMYfcLffzIworKkM+owdR+OVHRj0IKrd0byegJX
WQi9sT1BFDMz/PGhf5+DpGceFJ7heCTskNecAQyJMdLeKtkXy+h3x/0ByhK8OAgBQno9Aiw1xHMT
nrgjvJnSg1LMR0WjYy6HdULUbp+LgAdcKj4ItRsf3MDVuot9+h7isTdKg/ExMgFb9jNMk1QAS1m7
iL23+Dz8fGAcLyZcamo0lym59bNfyqq/LLgZcn6MaH8hRzY4RuM0CxyJDcmEbpMB61Ev2BcWctQT
3sKxvQcWoFOJSwiupLWziINjQbj9gz/7divKYWcuhWi4NcfNWUequd9vnCwrgkEdHCE2MsljynFI
YG8RiEGowwKI5kzjd31IdEywTROAnAgEPFd3Z8la4TsfsnVqDlqLJfXbXLz0XYblT4AkAx2cEKz/
Bw8T6foDa+TDBViN0vfTRKlQgoUzGJDtmkw9SYisXJueFxIqKltJVyhY1mHFn6h0KRapU6CoXUby
Oi+KehEvtb4em1yQNFIgPJO3LcHIMtEy962CrHRoX8oM+V/mJLW82j8GEL42nKdGdPbDecEsDkvB
yVx4arx5orruk0dGWxk1X3d1V4il42qB9X8P1lFNzD6+szA4JJz1/e4AoTuYbCKwQoquA//auohs
Ky2v3twzOwOpu5R8q5eUjI6aawNY1wkABuSBfSlEreYm4Yjls/A8cjoD7mW/b1H/DBjFbwurGKet
sWGBe5jK/lXAm9lJjWob0l0JD3ZSmV5ULyN2iQHWNZv+eoAzGz0T1cBsIyYFsQh1slQC9MWuFag+
eebT3UO6vMfNhqjgp3jt/uOASDZcI8ErctzA7GNCKYzTiXWoOKYtqwwnhfBv3o+yzJ9mcrEEzPUe
7mlkuxlteEP4+bnjY6/AMRma8ki1bwCD1MouGK+/Y1qB8SWKchWD6odHhhKFAz3yg06xpOdioFF/
RKGePYvMZoh62HGa/dBl8Kz5DuM/yjnZHnPUDa/dl2rp9HjNC1gFlSWGrEqr8fftndgpU4Jy00x3
KTjqpi0/zpjSUSBbqT7ASE4W1CSsxvPuZn9uBPl85bfSH9OEsorGVQhm5198NO0Zlgw3ZP8nndu6
Dpc67CYSTD0T/adhtP31WRE+2MDzUCwNZ/ezOEU1LFs6ZLEkh32FNtRYcY6aLEk8GmhoWnZqSivZ
jKm4dMO11f+ETXnQNEUSlTt/fuo/Ph2N3I5u8q8cCz8sbzK/DpN6F42QPnN/hvJ5OMFSjbwyf0nV
cQrTMq5h+2RIF8Yk/y7KXoWTr6TZAnIz7omwY7ozEL6IDNAxkkXtgL3ZqnT0S9IpO0o0rZUVln3w
Q5174Zs1An/C0tdAOw0+uF2lINfCIOMGojvtg8qvO0PUZkYS7M1pb5cp9ihPKsaaS5rTOC+9Zki/
TDILV2EJ6cBvmRPdL4j6JnS77YGpY65N8Hs/OxDw70RMDmmh45hC+odaX37y7s2nPdXs8roSPNP4
O0jM5xluqDep5PWktjnQrghxyNErn9hjgxmag5r6wqTBmXZrijsvfvUiOJwNJQjK7w2qQ47JJ5DZ
ivsV3WmS6fIJtAYMDqFP5WWLtMzZwaOQJwkUJTFhjzZGsp5ry8IU1AuVie2UDMunQBiiYtygoA5p
wavCvm+Pkq4mCz328wcwZ92EbEtI5p2eHB6xQo+pYkbvmYME3gsvQMi4FrxVvkphZXes8BKZg8fr
k5uFxV6N1ectSqe3a4S7scmvss0EmPriMp7/YhFdGRaLqWz9xpyjYWT5JNdQCbBEgLGP6TS3kA68
Spak0Jc1ZB6FvPGEzSLIx9BAbn6ytyFVzE0dhSeUHhrTT7ouMeXFm0UJnWZ7kQ75jWzg5yhcjFdn
2Greo2qssLvtbrpwyNeC4HuBQ4ieQkkDiuLRUm9T+tlITUtqtUVJL/jXeOQYC950JE4BhXrgzCj4
AxkQRzI0PjeOL7Yj1dRO1SqrFrhoWHvHbz2POmDlMmX2CQXNd9Ef2m1d4cwkaY178OVXSf9exh2v
+DK89Z50fKC2QU2SHBzHXNtzHtpwo6PBm15nA9tAFSqKtb1PoU1B9vwfXLs8U/Oil00kln/tV/Lb
HDNol9ds6d+tAISdYabjuHEcDygYgNKDKSl3fdj+v2S90jvcSqxxth4FLwj9/No0ly74FDMmmyNd
1xPJXzKkg6fwuSZS6suhPKUwGOUwvFB0XLwHLzgZvZPm3TQilHf9PySZWr3Qlg+uqxUdPGxQcYvj
si4dWi7OjN7Xbl7P8YC0fPuccixewkgb+EBPicFz45QUnvSkPyI+eC8XKOLBx1vR4eDQiCdVqSha
B7QHTbSXsBhk+/XhMBnr6cYq44AM8skW0bCj6FpU4fYFpxy/6Ev5tPgsUQh8SvIOv788qXo/Lart
CD6rTLilG86sH+1pI7SdJeNWuti9EOWbcO0yOHvgBa1tsqSeuGGmVaACE2RN4YjTQhCEWa1OH/0X
xf+kh91hFqPzbZ59uwh5r+df2zhtQsnzyd4nEqtQLSghlKbyww6PNDvy6fURohtcMTQROQUPA/aW
uaUOExpXMR2exg2/Hn2ET7CnW35H/RhjRNYclDG0o1S6xxvTTY5MPScSzArgLnv1zTLhJWMbIbph
hJEw7ygOkmccWXe00wygyL+XdOQe+cYhXpBW5q9Er8+7twKKXgfRgzVCjDCVTM+3kSUqCrvV3f+n
IGgponTky8T3PrHsPqgWocNZhEJxgu23gTzD+43ulDCeV/DMK3dHKKk1UknVLcRmSeeOodCC9uq4
MTG3d/JL6vbhdT9/KwGew0MvlASc62uVKjEOkp4UjVYPVMEztjAn7Gn6MbCcBHWNKUMsUMUtiC/z
0ZUEXgFPcWDdaZo5TX7xyh/YKzTAITgDxoN8WlTyobSPCHlDYMhKeyjUKX8f6pHa9i128+GDFpUZ
PKfuNE+t5zpdOqKHd/kxO5U0PACasovBk+U+oqUURNYsZnahaIXQiiA5q/Nn7gJSJY3m344vCzBg
UlrrHMTnG0UVVls1VfAYdmr5thOWltjsQqDVhKz53+saAs4FRSG5mreHHo1Z7naG4jrJeXDasH48
I31rDLoQ479C2TMDH+V7IvJ90udi0N4Z31JDF/07klGrzZ8c83LYtOSAg8G2i5nvOOW952jKSE+1
SBrjjaSmP9XanPK90DDsqkkfzq63PFwDz5H474F4kzcj62mgKv17AvzZ5ejMSrhQgBTKBstb0l+q
E3BEn0WZRTmfMZJ+MwlKC6+O3sEXQ6c40fZXoVzMBqUtycagCF58y4b2VjwfA1RGgm/nMP/ujkaa
A+Ph5jDNPyr6eaxAx08gs5qtd6Kmg6NgLiJjSnQsNTJnpIe6gzP1PqVoQPJFUcAICnZc7FqJw5vZ
kfIF0uvbZV8rDctKzXhmaPpWvbKypyWBLoExjaIdANyO3+2f2hsHgZeL6+T5TL25T0N+V0JMXrLJ
BexZT0g1pRdziIGEUaVw/vZCoIlFIVAGAFlG1IMyaDdBMo8LIrqAzJq98W7hRuoZYkA1T6uWK0Ov
dkuEootaz6KMA3GBxD0Z9VFWYlaYhYeKE+vGy+mxb+SDYNaLuSXH+EfdLoE0fjhnDWuAadwVJZCE
ZaU9JhfDz+Se0D9jIn4CH2QH8B476yEY0ZPvhAHY75CYZm6tLy6WCaIhyhByVl7UY3H7VHCqgc3f
546xKJbBWCfOth3POjU95eF4uFMigubHQJyhmiZLCKFOw0eWKyJ6b8XDIbVjCDz48kt52p9BvQfi
pmvIDwBfYKkzumT1mynmaaG5DSxAlVT2oi8nl6bHXKehZu0b+QFEt2a24q00udxUYocKYfr/gTPt
P2UH/kJQC+VSZS/iTb72nJO7AY8cZomH5JlIEMwLEQ7q8IiE1WEBKF9OnWtS64i6DLPlyDz2SKbG
enXK7vcf8USTzW4EobT0x/Qt51TY0Z8vqpOZcsPiFfqV2f/t+rmaWyUyXIcCMDOmJ35ucoYWrkCH
oYRsFan7WWoljfbB+Db7cJBK8AGh1PGN5ahZzrb15GJLMfIYEne6U8zpayS0vREB5QMF7IxamI5s
R8vI8N7EIymoDT9dO8t5oT0KtA7Bew8MXgjFnypuemmE0A09zTMt67qZlYsGDCIbr7L440VnLZfG
Y8NC57xsVRt0ypTD9nAokQrKZga4Kfh7QG+vdva4NOg2yhuHJuedKeLQPbh+uL3Y3jFGO2pMAldb
YmZaBA4EQJMR+IrbU2vrSddxZMEVnJTuRp2lmesRCAWMMIkJJ7j5BCKyAlGfN9qVURlOEFgua363
dCTd2v4354w7ShBn5Zj4tGi5eTVqR+1bPDeYinYbRMHwUA6I6QYQDMiAplGEhBKVxT2TrE+MpXTE
D8QrzEPbY9SOQ6NLgJNZJCp8sW4UTvGc3u1kJm7zZcrjmRt/u44BAs5IzLGX9ISUDG3LnBsoEN3F
pAGn4yyKvBLg3KgVr2v0xHt/YawngTPIp8JJfhOwekq19doTo9ORc6k3VjyQenbnhqPR1zH9SEoc
4rDN6oG6cYdLiPVWpm6ph9/KZ+NYY0wPywDSisvfn9JpQ9D9wnRUdAaxmxFSMSRqUt2lHKfvw0JP
wo3zZCEvqT9sFbylNSsBw01l5cRVu6yF3SSqHnrL01kC+uN2kG6dnEMvYsIuIyN+r1GUNKBO1WZZ
Z1wFiCbBdHEf9vjD19bRSQHRmExpFhWT5iauOygAnMZpyK96hH1yOhdabOA3hpH7fk4QJxDtZ88d
pBl85OOf3zgeBR8DA5Ls4RmtJeIIrJC0OPxbSFyteewh3AqjaBqVbdozxe53A7SvvSi4UAjYeZHu
zmRYY2+f/f9JIniq2BNTT7H4LtDcWeqM4hlQcnYLUusJ3ZatcIJXIQa4SFbJ86fNKJq2IgusQoNN
CYWyCopQjzv1bkY9nDJP8DnC+ndWa2AsML9/vj4q4GkVm4EELjf+KiXUEg6zmZbkc6lk5CVOGAyJ
8gSQ1C3xAlcJ0klIe3P9rSBsIV0tpibg/ecPa92kLx5hAouuPbveYWiC0AzeLAswnV0hf6cwkiFs
ooMRrbtp0YVohpDvqYJtnQWhyxLSSKafgZ66WsjRX8MoKPbh1PooBoXzdfPKXc2LqS5gk4M5ia6V
bGxU+INn0LJwkwpfIq/PgoOn702QJLg6Q6uUqPAtW5CjEyyDUDPaz9QPY+E36jZzxw6LOo/yF6cd
G+M3q0QvKriFbL1W7+p/vEl7z1qeYBcqOR+tBCo8p1zweWNZwEmM0w6oUHPXIJvS707h6wD2NBxc
F1slkg4168GWBsC7xIqYqAbjKYNyAAkDzaY4io2NTL2ViGiTBlCXzCryxF+9FfP+qll958VOlInD
KNJh6LD33FsV6zkpQR6kxIUA4jNuLNprHP7Tssyt7rqH+uEBcXBk/3bzCINog1d9seDYzSzAmHSS
QfWtuPcLOMEHc4hrp3l+5cxTstkSdO/KLMl8MZxYrBcrYt9pq0iPJGxxNyQtEA+H8CCnYmLI7abw
kZRvG73NXTJTdsVv/yai5rUHUnxDkdx1hJ/jKHKKRDj66yXAPQ0/yx/cWFnVszxO/0OJ7/mHf1Fu
b8JZE3mVOqAYwfvR1Ls6QA/xfi6G+jvb6MvSGx+bCrSgikO19IGNtxVFNkSs8Q5pzR+s6UVUaLb2
x5N6S2saKzkacWuW/gAr8Z8LR3vZcScIe5DvtEUoWCnaEkqtYKwNHXNCOJzws7W+ME/5AyBAes44
Qf7T+Tky5D/tNUGoklPrMgrs9626J/XC7Z+HZx3I1be0iYQyArXklBF+85Cxk0QaiXDQLXi1T8wR
X3HUjd/HttD9ynRQrxj/1jd/9f4QpPyxeJkGNROzJ1iMOL6VTato/X/rMS5H21rSHxv1m4mPce0c
lneW0ZxcAlWOHehgADcft43AAowK+KsJx+9Hgk+IXkEtUNm1vgA2+zgWMdtG1RpLD/R6/XHdEb4f
6m6dcvuc76a1mTnvRt0mFg7NdWPOqckTIxTDhxZ4B7LhW66/mzs/7n96tvlyAYEwOwS4oQiQ2ZSE
JtRUIki5RuvkJZwfJ8fkuYlACUpCVHLldZ7YVpBsS8m1hJlY56Sbj6CDRP4bK2q69Q0vOer2DzPR
xwn1Mug6WqM5PlT9zfdAhLuSbxAMdhEIi9YlcVPn+TL471INUJbMgAoaq+uU/WguBVH2ozTrt7dR
tRQw97O5kNjy3QvkT4D0/h2ZRp2BwxXRjRH3TRnADZS7FoRtEgN0sXdYZSzpkWvmNmymtHkKH1eh
mDgPmXxttwZTtKK6OFuwLLU/N0rioH+JKf30xY0/Z7iXd86F2by/AuCUQNltQrasd3XqI6PKVrln
79013/07IYkOYE/e9CozYGDUBk3df2OK6VEGRckoahU1A0cXi94Rd79/7/XzwxpsSRa01dw/YVv1
ekwS1jJHQpqv+2JoOYFJaSPYA3wBaows/m17281ya0HT5DI68sP8pMMuJPC15TT3pTiPPEVjDyzZ
60DL0ffUPZX0bcB2CXdlYUa6a+aOawXYmygJuyad/RTxQXABVi6gMaDQ166xzwBTpSifkpX4irvr
nN59niXXjb2RiQQDBe0NQTG2AU8ygNk8tEheHpzNGyUlJuua4QvSwnF6NwqyEbLwlzyxPYetIIGV
1vpiBFYJUkC4WNcweue7lqQklchqCiNP+rs0Za1Xn35bJuRN78S25HSL36x2LfqTAnbwmbJJSNaZ
rNz6sLveVxSrVvz2kyF/VjXMV9A2251K8+iFbWUXGQRu72/Ay1lyYnhD0URmc8bmHueQdXck64Rk
F+7PPd5UdhMaIArsYCGpnxcALlbG07H3B8SCxEkTC+I/LLxKFh1XByPJqWegZNf1MfjAYM6lLjjh
tIXqcnHy5F0WR/A3/i8p5IYQtURfketcsWUrz1spTdPIQi73K4ajWrdifZ/tWZR5cJO0z8Qzfeqc
dj8gxvTvUBEFfi1/zgCY43o4xs3/r+IFvHeEXvI7T1vqQ7I9mwy8WlcV/d327y18HxSis2Pc7UqQ
pfKhh64Xrhc4VPK3GD06wsU1He5ML662c76iHMBouPzTev3YbjpaNZmhGCYRBsC8qIYcnhaTBv6x
QClBmbTloALQQ39RsUjP90jnsBP3u9Q/99Zh88cekE2Y6W5HFxNj+//g6+LywDQ6C3A6kYlykMV7
Qf9lgG1An/ZCadM97H3vEGHMSY6dfq/52sbe0XMJ2nO4jJnEnWlKkFIpBk2/RlcR2JLJ+n4RbvgU
rgD5zGKgdgosphz1l5b13eMdkON8nOadPkltN5srAiTNfdvrxmM5cZbPwXU3ew2pcppLNjQHSpN5
AwX3Alydx86QC0yejoMRHf3n9k6Opc6dYSwR5zZP68Dkyjxgzbg361+YIQsWFXU8xDlni9zSmnt3
f732mgv1+BVkeBeDZVBa1+/9sPfx22+w57hzvbGg4Y3kCal4bAK4aZIyOmBJ7dNwrvEvcgXxABxd
ecHqq/B4YsH1bOtnqqIuKff0iVRh8vns4ecXWoLaRdFdZjQOv/Ji6xTN5eKrmrozua1ccJO/x0z7
aOzY5HjZSE5glbXZGkEWWLT9wuY47OfYcxOLoKK9AQIawf7rOWHTIL8ci9OQo4uBds/rCssjedBx
7iqXwoQz8363I1U8o9YAVjqe2CqHTMqT6t4Jo00du58xJyOeOX/ABLkN4nAju1D6d4zTDlNO7lf0
XPXdqVvXl5LRbcen+qH/1KubKnCJIGLmwBl+qxdx3bqyg+OjvxYk17TvKD7/H/zE5GwwYq29VF+/
enlCRmpQhMtLau/o45fEGOt+kEUzhVxS+GgPIifCR3ipEu5NVshBLv7rUCLYYarGARIxbtnZq2sV
GBttq0dOd+GYy6C0KrUg5/vCQb8qrrrNidi/91im6vEtCarDop2S169R64MuQkI9XlLRfl1MgN/k
CJW7TDJn2XwZtgneJSrm9cnRHXI72T0Z4kA88c+qmXvUAPqvrOacCtgbD8EyCzIc//9hovc8AFSX
FEVthwMBrS2kWWAVetR+eMgDjVtYel52iPw4Vm6RJR0W400ws+nZIbafcyPmvpZs7y7OQ5pB1PGR
eOSHixV5lISNtMP7wPn6u4rv3jo/QE2BsTHtdmxatojKEbMuMfzF6BL1xzZG1inyjrEIJLy3OkOK
Dfa+kd771U1mG9X/aMZafPc6nfTXcHHI6orwa83+eW1G6a36iiGPEvOPI1e+4XKMYToGRxKJrV3i
AWsTCxyXvgadBovvP9cX7vONab47utEoazG/Xf6GuMCFFRCG0AmV65clJ2sERlqlX53LQC/l93qX
aeP5BE1khFtG5RRs+gKu5BNxeCdx6QBdal6jomG1ug2FdHYRI+Lfqpt4399ROjaJ3I4AYH8evkyx
osh67J8z2mWsVQXwY5pfWaFYfbPR9xGWobFtztKXW1Ewf3srBQJgqcyFyzLIWMIXy8/kHkrsJxRS
BOKBGRCoGaZdZeBOhO5vow21OaxsSSeglrvI1/dlDW1jL+W46tMgLV6s0YVgTdCJos/lDaxwyya7
WCmbUUiQjQay7QqBKuHQTrWODaiUrLfnTs5AvUjtPWtytGU1lzK3KEmQx7FthUMBm2B0G4+2I8lr
Rtv1iUP7Xq1aPM2Ec+dqSRY7v5qcduwhhn+Dv2yYe+46XAe1nNs0fbVNnesS6B4acddUHNrd/iwF
lyFGA5Nfb0sAqqrdeRazva6UvScf6ry4jXDGexxBxkL/lpTTLUc3qMCzK54ExAlISAyZDupczH8f
BzcB/hUJ0BU0wir34Da2uIxD1uHAN2IBFcXJA4Tt6nXl1OqtZdXgdIzIBfN2hRZYu6DqSq6rIQUR
MhdkWKqSmPdxq/OtkRpfFuoGNV1awq+jfifEWrcKZJW/r7ayZPvTHKXeqCyNZur56kywsbOzbnFv
Gwq4YPqCWqoqmaLNfXK1e/VKlY8kU127QaeoGRSbR7m24qU0nkpcqBuU6QuAeI9nj9CxXs4G8YeR
xtROeLMvbgsOOjGXgyg6rXorl0kFjS3Hbtif91NHjz1cvYcmHBTQ/SxchVr+BNisyvytXONyqL/v
lWaSjdlOg9oGXMFgpsIBfb/VjGyPUjb0MpyGP0KI7blxIUZJexjyhi2/LNbD+/5kx53YvKGAI79s
CDccgQgMPbGn9UoWy941ZMqWaDWWyfKfJ70eCMH0WspipLTuflZl9BxoV5DVXYl9Kr7WOjST9C08
ys30lkGCd4ohQUYJ98YoIgHtJ3EWLPWjwCCZEWT7GnJ1t1wHrDQ4CGxQ1JwCMRBeFOlzaJ1Z2Ikr
CZjOM8BrssHSVCx8pT760Q0hRhNLFMh91qGjW0QIu09CIMrg9XYnYRQ+KNnOFqEuwLgt5KCXFEp9
sYpi1xeJdGYIHembsaVqdZJKndIQqo9KrVYOZfS4TvyhW7IL+a6QTcdEh5m85C2jr0xAzkpU7u2p
NowMjra51tIuLLnyLymm0pc0EVbbU/4bJIojVxLVSQeJyg3QwKdMkl18s5+IR77ABrSB623N0svS
U2YgQ88+IYDybSs3SpeRbJD48qFi4aarqqEjMQWuHOvvr3i9VAKU50Nvy+KxGq1ZC4yWWQmWC7bu
emwxgc8tHiQweTZzs/7BfIGGB87BuC8XLA93x8e0OOmmIe3autr96q2vrHMEr76yTVhx6f+R2cEx
AibUOrZ6Xg8h5nCFA8n6L5dRBPf2ODJpw3gy2y+fKX6JVsSk0o41cbUHI3+Pt4tz0Ao8oAGX4FOL
OzzYbQN9SkKQu4B9k5ghpG1uwIXSO3CU4UdCbVE9ZUG37L2mZdMNPzcYEf0ztpzXYU9o0BobSIdR
2SNhzVP1mW7lQwLMUZcKwd8g0XLU8+lM3BKNOTnZa+BANb5SQNiR5aYFhy/EDskzUNN7DDuYcOCL
lHzGhwNt+WurbALHJ6zrMtKFsDWHWTe4vWiq/zEusqhFeTprVOlmPm5OIECOqKr/i5/SPediDed1
+zp4lMavYNvrXYoqAt35iwY1PzYeipb/qh2QRuOfgRAMSFpdGI+dZ5gpEA7la48PSh/e6rRwpHd9
zdBBJ+FfklY3lo4j7M/nvCFmfFlls2YT/8rRz99cUO20Qk8sLnPcs1gX8PwVGYKnHTth5qBS4psw
J9sxR4eoHmbUt2CiCMX2k9ecJQaI4q+6/AqRp4P89YPW52kA6Dgo5tq9O/JufWoYbs1P7fgBkL2L
Odi1uR+JUay7PEoPz3t0LwbI5CwYwSXpikrGRoM+dWnrxXQx/+7Zs+vcZFRVtMSMntacQ9RQsGoY
pVPWdSG0frc1heTLUW0LuGGt16kUJp8C6MANjpS4s3vr0/71vt4iYLKdah8kdXQ6e0M3qGhdi4Vq
pMjpe3iSkN+ckGG6+njsEfY/KzO0gnOhnLHgOM3aG6y3NBI4Koyh+9xxaUQS08HYg89JZO6hAaiG
8uG737yL8YzXOk4RSTQb0KMHuxnlpiKgFW15ejnMKL5c0cN1aZVZ+xtq/wX1solVWCw3PeUq2t/K
wjmkVqEUsazD0P89oOzrT10GvEiRE4GbiyFn3N3gAAoLlhOkMMV3mtD6V2yvBcF2gc3yiESln0p+
WHqahP2MWZ6JHQ4RrSXG93yjE+ojAMhVZDBZegiwopnI9vIkL8+CgbeffINrkr/ztxyrTBZ+mQed
KVEWqCnlxfhCIgRHPR4R56EyCxNqcbPvNU02vroNamYCeVFgnP2Rp/syLArxX/acC/LOJT4VWiIH
elR5X3wLbrkTLiuKEUx/nGMvWNLYnarchaKxLGO5sGW1D+waiIZ4dTVaK0Fx0mkVZnhj2o3upWPO
+hM9d9FcRk2TGZ5GmIW4wUclk9vQYLvveI9DXMRzsZpK7HqFieDnSD7JuJ52OQC5kJGxXlsgo2yN
nV8RGX95OmoJ8JgMaC0gfO3sWl2AA4/Txr9NKdeImQbi8QZ49bAsu3/576Xe8dyYMGsHYzpWEr53
oUro2cqK8NlYpdgK7zbP3zYPQLrxmkaQcsB8twX0anXwVHXDnQgMA7Mf3nxM1RuWCdscbj85vtoA
Nydww6MaqgDYICNI9Z5yF2dRngHorDyF8lbBu4PnlEOpFq6+ddzAfKE7j6KqtJZn0RTtI6kVmAjV
txaKTxhRnY8J966lOM72gytu/Mc0MSwZWeJkDqY0Pi0wArN+rZsqWIJqrsVDhfG1o5VVsG3YS1Wb
oOcqN+I1r40wudnCAt1jBQak6ABrX15ZE3GmG3ur+s29R22gMAsXJfibivNK/XNwh+ZbSWeyu4RS
wxLPmIUzVfevh4mZv4E2CMbT34IbaRqeqshyul4rkeqk0irdq8Y80Uk+5KFHjJpjEtjgD95N53+o
cJg8cII/4v/LwZDyzg712CUSkbrj8Gg1Uc6gHGIvmmpO7UNL+MKjEqJNkE//y96Z99VnpX13VJ1D
qNeABFTQezNFW3MHnoP4VXDeZZiTVSkY05ouZoox5PiKLNhPg3f1q99Wi/Y+FHUKvYYVpXuUqnKc
5EPKthx96S3mk/5YlwsybefBau/CpR7TSQxq1ZOU+RZPdT7RjnHaYbOMqEoXf8ac/kFI/d4JG5bR
Wzw5Snwhd3bjLFzZzpWZcd3Zj3cEf4sfCrdUDtgFdyo7199AoJjHyNUHWbtWX2QMqFpXF3Wn9NIJ
FEYvQBdV85rBE64sI+E8ytkJRt/fp/h26eam3Lnh+Wj/v0Q5jV3Np+aVCMJrGE0Ik9A+XSG5WFS0
GEvyRuDhSkUb/CTZ+z195lQwUbmL0UiN+Wr+hMZTFkOKKZfsk1B+Cvjbg2cGP6lUFtiCZQRyeVZH
v+ro04pMYxnPWLHDkuxOceLox0coRjfdPueT7Zt2le3zfw4ogcBoZJs+Y/f/BikG4ezuVMThnC8h
9KmiP+uewkORjZS5q6N2jolYxWJBD6cSfIUSP8Ifb/VJcbINiVJlyQNwU1cyPQLXHgQ6dJivU35n
JzatFTTicayVXZhEYSNSUUj7axF0vj0SRvvafTx4c8z78u5DQpxXS7aiGsKNDZ6KH2Bv+Jg90nwY
dL0Vyap/lkf05vKWStsHUDV+4nMnKiikj6e5W/BoY6O2nvYMe0FugxbPSEzE51juZB+7qRyoKiL0
QP63U86pnG+0il48HO2P2g5TQamZ40tvN3aEp/ixIQCOa266teKee261590dxJztc3d7i9eyalTm
PCF3uEpyDS84f3mDVLalMSoV/a4PImn4l37oYbTtKT6Mk/qsD6QYYYvis72kwlE7fAGreWsOBi/v
xBx6VfCyb8cpnlK3Ixt61Kam121lPqcRr9cgXU29IxenU2BpVLT/TQ1As0RVgPsztiyO7Kw55drB
PYdFsvu6zIBaBz/5oQClrD5d9xvb2TEL1B9jV6ihlxmszQ+SbGqVxJIKb03SHxmXGopA5KGiwMEH
5kCwjOUsbFLqKSk79721GKPYwbSy35RkAsYNDlwN/IIFReeN5BcR9jHpawkusYeYswg38YNwNyX1
Uoqweclbs/r4t13Qefi/xEU4tfA25usqR8aM5I4f7kSnsh06Moyc57aIUvhFJbDAaRnn64XGomir
tc1e3ZHOTPDP1dJeItzepLwL2ZO6vVVhDRoh5Y95BSMj46GwmUDGe08XxZN9GB5zDYyQX0ZsIzAU
UVHNwn2pyhIzdm1DWXtuiEHFh0ISgmYzYzotfRy6SaCqzdfxEGDAxujnBywasXO8Gpb1amuH2pWm
+mKk7BkuB1TlZnD05qgjwj5n6PRYa435cBGuXIquxdGje/dpRcbjDasECoQu8cXQ2oIyHGTtyYdY
QIjTiT0R4/TIX68loDDqRJ+0nWa+nSvL3pZJ5CTEJqnGSgdb6bcEpVxoM/M4lqh9DegNtk/NN0xe
uspY4UjoTktND2lDVdkKtySNJci9szAOjHSzmbrK9nsI1qhu6qC5AyJfkQiMD2IpZRktZ3Jq7pJ0
a+aXEjWxfurU4gWiY/fqKrnpuShRJPasWbIA7n4kOa9ltiEPWR70hTyqmCLmfsDYFpZCA2icavZO
kl5ztTzE63Q7GBBfrLExmMlXH5cZdHTE8uxM/El3Jse7/dKq6Hd2VMtb4Gdg+fRYCl5gStzwyXLX
r3qOQckXaAIG4eE9JXVgJ3EdTP2JxuIq4c9egjU8vOA2+kMdvlvM5ucGrKanpyFScP3fGHkXiRUQ
Ga+IGX/w/4qakeVWNSL9/E69iUawTdgswRTLQZwkGHio9caTIHgi+9Ya4nYSF7V0zIwr1cBAuQwo
rqhYPk4alYSO4qjIrQssD5mQZ3DqEaejeJ2q9D/u5FDi1jYrtb+w39fS25hmDm9D6KEC9N5p5BP1
M+E2rmNtlnCP6A5yo5Am7x8g0w/GEY8lhhLQqlUW/r7wFauhJR9KpY6Vr7ZZidjv/hjCcFSqJvZS
Kr79uZzPtyqo/Tsd24/OKO54LeN3c06tNNQo36mK9+yeWxbfz68agUshLHiYvSJfe7BmxiHSaZEX
mLxDqhOdJ5202pIKwZNnr15ECGbjgIa2yKdLXkokAdge0gNSwstrG8fT2Lw+1c8fIMPQQpB3HWBg
70TvC+6aDgLK1S8mm0jq3UHNiwx3gKq25mGPe63HYV+hGfxxVND86BYbDTNY8Y/KoWuoZ2CPURc7
S69ZMyaFpkT7cdBjZczv0+81IpXfbPXNQb89LKNfeO5MIK54FXO/mBBIcWs5r3SshFLV/2JNeJIl
/IXjNegDvYhdX3zop8hsi4MZTGbmRemFmdzKfZqFFcc+kwRUEU8FPUvpMoPQ4ZBJhp1P+Iaq7ces
o99hSlTFqFf+YMGggoi50Ku8mQAeNXoSecIlwQDL7ojdvHMqJGq+FJudUc9gT0+XSKSLf8ynqyNq
pkLfXp9dTD2DgrKukl1lENPFa9YC3e+x7W6reGf4WD/xJOz2LIfu0irowgvXmGkZMx1i9P8jhyP8
bGklEpQvBnwaMX1SYhl5G9/UTYCIKb40klONbhbwsk+bA0onIU56388A5Ri1sDjdIqxg9bGfn+WJ
wnbq//OmERCIUsbk+Zcb4ZKVQUf/aNQjAzU98JE8ft4s56rUWgcHFW5HEovqkJNlufDmBlGUojn6
X2jDMsvq8ojX84mJcp5hORn/TXEQy30lNUz0vUyHa6RiHO2YhA4K/IvSy7mVcCKH8ADZGYT2ouQ9
HXdGEg+ExyFXk7FJaaTElZBWJ/edMvuBVtb5nLgt89z6Oit+PBKv7NKChrc49zGaHxuOeQYO1Byw
Hsx4heoS3sOGXOJBFKJhPU9Cc1W8jFItdHhr0Ri8B5ZUs3OZ2TxseeMJ9MbweIhkWUz5LA1T4R0C
msUhMbfxoflfkI/j8pKgdVF4le2/wvjebVuJMPXVOjhq3aojPGHkRDbLNKUGBBkTYaoJwVn8Twns
9+8ng6a50zx7lVAHg1ACt8UfIglEybtV+yC317epUZkjRDHCFBF85G9ALIUPAgRm9zoutt/Qqhjx
lJoUpNvxQdjDpIYAStHD6L//fr8wHGmchiNPR4/XjpW4ylNUq8lqfIlCKVJpELgYWi7pbmFtvc3N
sXg0WdaLM06bz/kpuoD6/Slp3H8/Foqd0rN47hsWFkHWgC5eKAVQl2mP3/acVUttWi4mXGQrcWhQ
oH/c8GOIjJaTFGBpYTOndUhzhHJfwboQ5E8WIw8iWKimunZbOW2T8fvQ88SapLR1KHRbPOfj8wWF
VRDgs+b2dn+kea3D+eFZisp7n6YsOJe0suOzypvzYS+BKZJT+929afSsQ63DB+OsyaJD3tm/4ky3
8035t/6oJ0FWHLWnbmdg/pDr7SvgOkIQnZyEQFfzOU6xYhr3BeMS3cO929SBLZ5FEwj1Wz1I8zHA
fcD73wGEzKOkPf94gvTV/lZy2ILzAc6V9PWYhGQvWhjV/z4RbTm5rE1oQvln3fjPaHx5+wYiKKwa
YJGcTgV784PzjdXIeDGbGIeRVdZDpSZqeOXNJcfysa5E4wxnfb/LCLzvhwkPuVqEUJtQBkydhh8J
gK9NcVIudPCVDfDLJvbVurVuMpG/f50ICJLl+UJxgx2cShD1Gu1LzQfBIfgntVbYXcDCne6gRa+Z
3UnBS4nCvs0OZ3RIf/lVtVlEAvCE7vQpZkgqnKfuhllSLWI2/ny+xpA2SJbGGxlZrHwUPd6uovqP
8rFuHC2Gif5DN8CnH8PlhB1q0m6MHLxJLvvKofDqkyX9Cmxiw34r23cjWxBNAPsb1NqGz8orFwh8
Uhrb5uHjOvZCXqwiSqF5y+qagn3nb0TCHPGa0nLcf7q41rZ2J0vQoI35vVpwUVJki9XgQ6xuQdFv
Xojkwh9Jb4PgjspmL1jcmIn7rK8XhUwhdG8udH+Qo1iNb5DAuwEJPoCYxJjA2CHv+hcXZcmHtPs1
boC/8J8ORYyRLG2rcoZII6poGjJDhwHwn/sLtcZqCFQE9vyD9ifXWWmdcMmxvRSKn6vI5Cu4/PIq
Lea1rzjXhWucyCYtk0srjlIn5cJONZzkl7VBHxQxGWvHxAJtrv0bhnK30YYjCh/OqSu+dRMjTl7v
Ev4UTLVpf4JvM26+8Q0o71lOvA9OHdGQtiWHJwVK1PaZfLhp2R3cm+xWZqJhyn6s78cxrOgECiZq
ZTAE5ooGWmSf8kgGabICBt8StjhCUivsa2yLU6V63jlSTZR43xMTBJJuJMW+9ucEdk9dG0EaXY0r
6c/1b2sUuYPaP8M5flwxWD16YmyePUtR3uwb/pmA0S0OjG3qmwo+yXVfyHzI9gn1c+DX9N3rpuE6
wCFW0BGOczWLGqEi2kHSS7FuXSLnOhCG8HcMOpl1hW8vrbguSkapfV4v9ZOmtoSueS6aYG2/HCkw
k60o7uuQXfiMBFwAiSdKMIQaQGmsz8RCVew5oNcMblarxIOfh/1WZd86gULnRwDnyYMMHZZSB1YJ
T6gsvJjL+9WGzmULAAHnkgRttAtEmYFQDMxkuhF7rZc9TwOrsXHuqQQq0VUyZxeSfMFZb9IJN8yc
LBVua0VFbGpL52wQ/vOt71yEOsMgCf3MronFV3km0swblXMI77NP6DeNbjCkIoTFjaBOYIbKlJG7
tkNCbCQGEAKgMW5JDu5vw+myNk0jmGzSRLWGgkJFVpW8QBvQb4WP7OeI7bXimF2eNyeJPgFI9JoX
RxwU5NwRA05RWmQwF0YMtumJX+oHB2xRMusvYCMuPfqCS3FNwu9DDyuDeHcPesTg1YrKhhCfFwl+
IbTcnvZbADtaNRf54rnpj5GO+SjoacPl5bFnNk51mjuuF3PHpxpcQRdob6/Yw4uOirtBIKM1g9m+
0chxorqZQzg1dbW859XHaWg3JEE1Zyz1l0eNa/0BX5EJi/bH9Iv9rdFIQzwRcqbgMY5M88ltOxXM
81ZwENTSmGK0qDFJ2/PacYc7suL1c+7aMd8I7HUF/Zi2OCBW2kCkuGCMiEAyihq3UvCC7kKHBCns
HwHfqpoyo9FdyJZMAnvEyjIezi/UZ185jJUX7ouHOEWScpejiIryMa2cmRSANsKuOhTdO5XhntTq
PfbP3PVb1mpFQKNz3nO4pdnco7ILyK8mLFOwBDoqyzYcMrqjvk75Zm3dCMn2ien1srg9Nu74StvM
gcxzPX6tsWb9xpoueO7zVZBJRpk8FVhPslEEEJLwflQKOheE8aSXATglbbSrJEv4poGWQjONz37e
SmNBb7WtzxO2XnlRnDvzlaQ8d0M90mD0vrLy3k/lBmY0oMxnssRThCcFH76JBgdtSuHpDY3FktCs
IM+2Ewj+UwhGohsuaZWV5s9q6iZqLpbU1aLJUsQ5C40HGatlzDC3IrWF5VNEDQTfMCjcWv++vumz
MsguEZ+grTqZlCEgp98wwAyFwtA7peqS25dxL9tYb1meXPsSwjJ1mliAs4P6ru40gUI7smsp+A0u
EwNP6+8+/U9ZD8PF5lGPBNoXZppTChhVGBi4no5zNXl5td0bUb1QubbTZ7U0TIKaWUMKigZnXEJA
QseHaT8wI3KBVQ2pRenNVA24elekwWkDc9+Hkc17/vDLlYHXvhWPUvl/joiwZFXDYKYOPDGkgIC2
S3+6ulMHo+wzYRIgPQ48t0Z/T/vPm6DkvsYXTkUkcKjtt9ZDQdkuefef3Zww2nQZE8DIRiFIS4Ec
CUpsUlMp2tfA4zqSLJ/cNNG+6SsJSiXPOoZJBxxkKrFkoAqM/o5lO9j5EeWL1+dg8RZnffuxmwRo
dtUXMWsJltbrjbZ5rxHRgLxMoQPQeqXYW+RoLPPZ4NaZe4C69LAXCb9GiL4apdM9XXkBVBWkbwn9
5Ywj+lj/TzbNUkFXrSSN+CBGdgMiq0ALMrMWf1kIg8uPqWG1xOKsH05SjSqGdG8umy2F2toQbZe8
e/J1woyg6asZzFg6IL4yGTHBdu+zjZEt+7h3vvCs60wzXq9xsra/8eOgONeBDLBC8BJ6oRVF4UoY
zcTKgi0xBII6ULGOyduEQaTMHSKI6FwL79S5sBc1XyAi1txqIyowayjY6Xnhuukxkpg3AZcEweiW
7gLqv51u0rxk+KsiT9hjrLPwvlXJO3PYaEbKMXFrKDeRzU32WLGgOTcqoIbUytWJhg7vRYuUt4CV
Sd0jJf3z1Wxe7L47jkd3rQs0HtrNhAuv4BnNiSjKRWB9s6blm2wTOFJ57Rmd3baKIfyQGyWeSpmd
1rZUD9M3UvdfbTeUNGopVKMJTLBVax0j0exaPPkzDapIGPbDewREOVGibT+7tG7l1WP8BXgscdNS
1AuHL2ByJzoUcrMNM1J/WFDjst7wYQ0mNvEnCOtnpM4A15EWovqHfNpwHC+u8u9agZfr5hieuAaU
GBfj+cP4LLcciDB6M2dCFoe4lF1WMYsIpTA/G4grsLLC1VFyN87jW2Vq7mI/u6+czi6psFKpFIFx
NaYFbv3c9vPwFy1/LsXYRzGJCpag3WsrSgiveLa4u606EjmoHJdYF0ryxTVtBG6GHPTAOTbVnfEF
VEtwVg3Vc3yvlOrWu2hmyIyG8MDk/kBcrTIXpAMIzNewj3+LmJdqUHYGIRwHua+kqdjmgiNkLKUP
G7PzeeqBYr4xrgn6D+R0rhIq8dvU7Tk8qti/+1WWW47Rqfs3gHBoGGNpaabEvtdz2Bj6nvbNXeRR
GZel4XCQ6lwsxbp8q+udfbof+2tY5hc3NSNNND1pzP5ZjaEqZ1LaN2GxPeDxdM53TXQNxdpfjYMU
UtwrLFVmpq09ecAw6M5k5AgXN0r6aWTZI01clY/4QCpxSQek5PukpmJFiR+pS+5aH28JgeAmVhUQ
CdkZjipBbh75Cmlqvcq4bPOKTb1dwv0CuImbAL0lzljPefXKJZUt9m/dvyW8Gmc8YJb7PtvwQn8z
lhwKaKq5AG3Amac/QjE/g8s3bTTR9ruOrwo/DN3JmJhEBt9c0EMy3j6ABljhkNALIXk5D590Cx36
dANV31JThh2zbaRxEpaSBgb0GZBJ0FjII0Zj2m5RgXWSKDlmEphX3FhQLxiJA3zP0NKDCoTd2vaz
pSOOqdQVv1S+NjwyNI9OrvYiYVIAton0ko/adXDohgX+saREODafegn4slPor1ufYi1ABIu0vzWU
hOEfCfiv4hHrJnRN7N0BjUMwqGtaHpIKZFdGECX/bjLDx3WLvehd1T2al0g58d+VHtHiWo2rGW6b
FSBeEzQANIBhjFkBEJSog6FjxVKGKshfwPM28QQOIPgoSaqourNZV+dwWcK90xS041F4hKyWUiQm
gKuxbV8aJVHaY+1wMG3qGarmFtbKPeTkTIcEcknRRfZYmQ1iryvtxwzLxtGXgVaZbxi1VcSQ/lQd
Dxp1KyydrxfdOKg+1OFquZQEWQRSMMRjuy6EjOhcG/mEkER5xUuaj4kUIeYnKZZCrJDLVisbCkIL
Lrhzo+KGdIb9k+xyPufmbo9KYEelk2UgcJZcJDpps9vIU3tZWQtkURSUWFFfv8BY3iNuLrdijsnt
z7HJf7EvGQ745dKfEgqFrEf4pv+z3G6i77DzPyESMiirhXe5VsfslepsAkWt5qiIEf5Qwy8bEnVZ
rg0kZ29ZNqW3K62OHttEE/oIweni4tWnaytmutAUxBZQKCF99hhXnD/hs7nguiTCUqG/gLMw9Tam
L24CZ7jWZZKMxWqqzqHu9YMbEGrbecVecEPV/K3XMk6ZpM6K5btFEjMlCYBgH7nw/PBFbQKVIA2Z
Dp1T8b4QwGVqy+xFEC1863JWhyWtlBiyfQwxAsPgt2RbJHxhfiv3/dduNvjCgQw6vTkqXb0Sgw6w
sSoJ3RAKPbAfZFpJ2AcBOWsInO5+p9DfSiq2VDVCAIZLb065vf5rep1oj7yXVNot0T8I1thRX6KQ
JHHTRZgXRx9t16M9PO3vi5dUg1GtJLLZZGZ2Mf+Ta3K8magtW/hrHEvjt9CMjYCYMxuYGNooAMJy
YqTFAVNKkieWns7KKKWjja6t7TtNDZNc2FyXtKFbeZH9Rjso6Oq2IeNrYb+No7l+YNI+f3etRxdm
dIyyUaw5qEE4pZT+FYJkMlUyEvKvJou7fYUxl6BGVgKaLeSRhW8SHVULDG7VnxZ+eho+uKLf8Pqq
2ZB3x1QfAMyjfHR+VfSTAMDgupUIejktFAPpVk9ep0howHkU0GIwlD7VyH4UmMpUBXwQbb/LCdgK
xoUXfnBWs+Is+qkqLDtJLQClAisPBoy/k7mEmS8AktxZw8QCw+Ya8nfL+XyGZosqgOpJ+y13YIto
ov1tUut9cnmPbAxUMqDdGCGwOm24xgwV0pGH9WeXBFxsritecEFHJjAd1Ex66D/t67N0wFmhm/Jp
yNzLooOvmuJ2kerfTM6q6xiFFu3lan89F0275OVONYH8TJbMhLjy0wb2hHb9594qRmwL4X4XlJQP
ZTSHuqyJyxj/tDwxtodesMYDuM/j8kfI5gNjN5agU7WvCcpnxAsZFqVDkrAx8/32MOpYCZFhf3N7
15RqLVHVilNLrphPdRizFsCezYWFrPbH8xN+rs77ce7IuJre7i0JxlyH70ANpFlodAlwp84pL1tv
DHX4nDAjjGzWvmISoqJjKvGwvJk7rb2fu1WcQgcyAUBns3uQ9j2a7j0iDCM1sh2vhGAVbMrpW9O0
0cJ+MmE3qxUz7fCVsciKTKc21gLmC8lBBjYcmB95XvKdKimna5McFvQEcXD8ZccjIbRshZtKwfJZ
93QBTFdbyf42xFT6e3IExnOPKJ8kBDLns4PdNXpSuo+9BMsY+fl5/GkwIpL5vUzWajaKSB4ecus5
ZnwKgz/tS0R8NlRFXdFvAXWDAfhAqQRP7Oese9qNwZwkPPGP7TG0x8CQ6cRf/S+CL0vmvVCYonoG
WZZoI9QVpBpl3GkHV885fHSw8X5Tmt9XqUOloftIEXm64O553Jgd22HzVvkRZjhF2YxFx+xXfYBR
IMjwG1qNSi8NQbNimfbqUWBq4lBznA22c7lSNssTnXsIoITQlPBtjik4n5a88GfNC7h9kSPDTXj+
h/CXvncRGRmOYxNlFQRRdnVRCKJOP6AH2fILyyFuDygfNW51Q9W3IuQLiItjuUkCbwbi9XaCkr0H
L5C8/tm9o7QXAkw+KMoepYIztBXlV9i+8WdjHHhY5yug8Ikl+eOS83l7xPgowQ7PhiJRAQ2edlz/
UzsnlhB9aTd34a1GbeIcHyFftCJ+6PULOQDYUOfWOQWDVAzx7sfJ9EJW/f99Ms0uHULDWwrzh6X3
RlfWQl7Y9Z/lqgbHaPtWHc3t7eQVZYz33ZkHWUCXfCb62zToSxEos2dtfEJsWqAGM56ICPcyl8hV
d3BCatjxrzZOJ0TWBlGIKhl0bbNJKDrtkExL/SvsxnjQT4GVyAgLA3n63hJS26EG2uhqmp3F/35i
RTkTdFxc4Xyo3W6PAsoWqOmt5/tAoei6PmkDtBMNEOzyXlFLNpnfcA4IIv0uFrfYJLPdCFnV3ZMs
a5VkQeszuv3kbeJ0w/ilGD6Vmcf+7/GcEVeUu4PAMoVfhuH8oUaSud9w/P9LmYlSM1/ZhL6xF3fr
zl6DT/pl69L/UTItsc7PKKialU+meivVZyJclKLc20U0gvPL6DJra+g/gkPZQEI6QO7k2PrT99ti
2hiDD+SvsPsg+5C8LSlzQDO9XCMbwlm9TOufcHqRykzz//gVU3E3j71vPg94IwdnqTwRj6ao3Qis
OIqwl7KEW77lkWPH8U+/eLwSuC2MiLDFZ2uAwqzrNODMEw6cA7fDw+ZaHC4oEY0UEQj75h6nx229
FxVIpXpNZUxuxFDYOjHVXqrxvXsgXi86zUv5umX0aWIJr/4mnmrlS+MuJA1VRDW9CxPbvRlvKLcj
LIPzPoWqZZEliwxBVxT3wY6Kl5hAMKuIcZ42qHZdHz3sNrovuvmU7C2nWEied5Vs8wvAQ/Df/M2N
iY7VTPfFBnIlGe6f1QuG4c1oaaj9thzrpJXB185V9JEeu0Hd9X64wIpPS/l2y4owN392oOJyh+8n
zdKU6kYXSaMFiPq6cOg0KX87ViTCpc/qFsk6efupOciUDAXgeL8CfATMJLpUjT6vColi1nGx9zHY
Hn16uXvNVKrEDhXxynJxy8vgRbRdsa9HgTGKNuncx7uWUxL80VV48kG0yXJ2i6wSzUYHBJXn9pzm
rEw90sKQYWmOz1OPyToxZJrYz+smIMid5gwLvhierjI8xCR6+4gbVzcttsvnALGvzTAkpSoR6AdR
/N0cla2wekmAgUG12wiy/jrPQ9Av51NKzM+54pS98SXWAo60nB0xlCl+MhRyS5xMCZ872ZHfd6jP
1wxW9Ef6Bu+DzCLF5XFIuCRdj5ZOhr5ZAmC4s4Kf+0rKtojwgLHKUQUUgJIjQACOc5oPNOohH9MT
dL6m1KU8C9xiwUR9JeijgwUgXtY2lFQL10+3IfXFRQZJlwXSAM/8U9kYed0ZXe1SNwRrWZ6Xx4P+
cVgAjv5QJ/Q4j5UuWaGA/+Pd/P6GwYkM18xCtpcB9SjkxD2V7XNP4hVfgJUmreVg/QopTglzdXIa
0YuPCdaYba9oDmWb8gipV2hSnGYURXg2hcsnRNFG0px0xSpmH/YzzK4mn0qvzZlJt7KrGFl4Np+/
GABDglw3TpQdSfkZx0AS+tJuctD2o32AyzIb3WIM5jMtILt/PMdINS2onUPiPtQHhaxp8y4CpdcV
mFa5YuZbPKduRmYyGbfobsQSvgoO+wn9CMTC9e6aXAuPYVEQ5sg0rqMPiAaoY8BGLTEl1Qz8DvnJ
AgwjZmSw4c631TTBtpuFE5I4OiU1iXh2MGgDHAOzdomAJRClKYX0vNDR9BwjN441O1K6RzwVYPIv
4fF7jlVKt2LmiX2c+Uo8zFrCfaj/2CBSYJO3WHqT6PRXMEOaZC6d+9jwwAtmig9ot+GwaiumKLog
pPqh8cJTM7fChdAq06OFKb0d+l6U7wtdMzwr01pLPxSSlHMjjuZMtZJux6lVMBTumNGoH+eIoH+y
63IFtAvRUVeLIdWYA2tFLUZcrAMlAZJ7Cfp+qrctyeP4liX8UbG6t/XIobhbqSYjt/qRK7pzBssv
lK8NYaLrE0ywgFNDfeV1ONBillwBVNoyp0raWs/K76GBUtKOGRVoB11cPsKDR4G7sFDeQCqYeYk2
fpWrx55CuOhqKxcGpiJcxLX5YhVCt6c+g9bV7bzVUXw+COWa0Qr0uPnGzwi/ba3WMH074MGyjH5W
YFsTCDf/+Ccqdhu00zz/vE/JKJTGg3bkIjHs9sWGU3ohdizNQ1+y9gX9dJB9LAcLELlRiW9VTkvP
/niZAanL3fdEcqbysm7ONoNSM59cTIdTS8dRDWTLzOLEkL+IoYCkDTX5EGTPlgZAqLEEWIOw1q33
Cp4NrwImapxttlyPFWKmobAykitDXfcPRWZtTaBijl8CghLJtxBfHLGu5c4r/BVn8XhAudMoGMfr
cgeZ8kq3sVzV94wGFsIFaMZm8p+N8uHCCuOBa3ThGxqCbG3r794zGFOrlWV13hiCczWdfrMobTww
BAyOh4IJbsMxJ33lV+q9ekxH1/TCVvZQetnSXHWp8uLzZM5mqic4jx+EKy4pUNkqJliUn6ny3/cR
XyPZcNzptqBHb/JBcn8RWW15FDVdzWWbKjzfDgwRSQ5z+ZGrps1I2HtXM+F5gIenaR6mZ9fz5a9B
bliOU6VBCdIMWq3xb6pDVqbUOubg65+AqUrB0YzkdmMDgRO/7/eVhTKHpWOUvp8ZErKlHRGP57YP
lDkl+YArLrcfUKGddIE9JbvCpMV1yvp0DlAb8JpwVY3Pm5cI9hOYVAOsdn8vV31PuPa7TIad7lUO
p8qsccjBiv8s+k7HNZl/CVWbLwuCZn5WD0aoOG4lSnuk1G7frkiy0jH7kH8x5uzdhoF9IC8IO5cu
0G/VzH3vaJaUELCU8/cs7rvCyPmoQxvaouIhdsPgPP3fZk2nTSOcC7c2VImp6ql4gz0G+543dLra
4QO2amkL3aluFNjBCQlEqDTkqHZBxFOgIfo68yEGG4WKbaa9juallsDg6cIV9pqI9rXDROVq1alK
MCX9iQ4a1Of7uExn66OibUt1ntMEsuZ/Lf6m22xbik0U70s38Sgw/KZ0frmlG2Alz6Nw3nktul/d
3Z8gZ1NYr5e09sDfCwgCWMzvWlBkZQKcqhtvEVE5P5/W9nH7XgkGekjcmch9WXl4ySb6QnrY9qI7
BnWIaD+AuqQguq+z7ZFXitCYJDnt6Ldg4ZIoM90vkjWA6buU1pri4JCV9Z4iagiqxyFBrtyUWNQg
jByb71z10TG5yGz6GN40sxC+46HhLKmtkREBYIo7AhRPBqluELMCW4V8L3UoduCAPTF+NhH9l5WG
+9ZLwiV1j+BTsheBiPFYmNWArHlKBjxK9I778vv4xyhcRcc1ZsTCedb+0CUhPcXCuCE1cyn/1ur8
kbo3A/mSbi0slO6gVlx5G/QXHPkZItZJibP5gzQ1b/AB3OwdORHA5iNLAQvMDvgDzGzIKhYqZtBs
7nk5Jf9D+NZXtpeLTsy5bGZVYMyiScvlgL9/fNk74DfJ1w+3lsF7SxqlkuD4YxgiyG48IR9XuDfp
pYHEBDliVx4qTe6q+Vn4a0aTvGcDq1lSuu7WpNAZVr77eK+0xcK3D07WwTx+Qem03BMWtYgsPjHR
AkHG2gSpU+R8I4KoKZRqQ4aCTxjd2L+xN2cbQxL48X2k466CeIVS6ZMnnkJdvNnI738EOT85UXWe
CrrqI5/CuzU2HaZnxs0GzPky7cVV1cBOydBz6BWExLl9rAvYxu4peNFbsZsDk5EIXi5abkylLjPG
qaBcdMNXZzBmWietkK/rR12x30TOovKa8iZS8SGgxsbXhWYnxBqFHHUb4dqW0mt5tUE1curdpO3x
QySFlTCOd1idnOMuKvLBibNPl9wyGCZsU6HezezAl0hSEa3QaSujt+IOc391EQ47x9Yr+7bbG0uY
7X7OSOMKmJUQnlmoFnNkno0cR7WGHcxPgqweY7S6V2CFcKTdbIYocsb2uS26IjNYng7X3bA55YUQ
kftNVdVQXgfF7AAhc1097ygLSabLXiElTvS293Hbg4Nr9Cn5wtA7ygqn15QLyt397fDrR8p1Boqw
BsNOhj2u026fvvNS2HjuttuRw6aAqjhm+fkFzJ4otWelJDUZT60nXo/sZMARIpDXWeAheMh+xm4e
rstZVbVVwNXJcUgldmVsbjxr6V2tTwq/gxuUbc+L6eAlitExedi08fS/DIswP/fTNx26+mEM/OuG
1qno8TWw3Gc1mqlsQsRXZ9mbjYgQmHe/kDXAYrRwJUF0NgSGCIg5/s8D/5C1VUHJzVzownKw74/1
XUNj/tC5epWENLbIkRrzEJG9Qf7ybGdeJUpCgizC8+iBa+N0Kzs4EnSHxAobNQAFHhJUIU8Li0aL
4bCVGxEClokBLWy2alMPBotfCNUBcxssMyPVzhPKAwXOuK7DLcpOVfkMR28n74Tr3BGn9qgo+eUe
4l7CMCuouBAGAqPBEb5tWcR36zFN+2ixZBUIIbIn6GP/HtPSByRT3G2dOzu7Dfmmw3rDDokP6OMj
d43l0yi7RwlUdgN+ykegYyuhlmINQnw/7v9LNb/Qiclh9Hs7Xx+Kmm3nixM8GH/ygPfQhcYdrqaQ
C/fDRzehi99AYluB0J3mGi+XZ2eerL4lxFPZQ8v+Ryv0JgijrV+rsWj+KRIdTtaDFSG27b07EFzM
3pl+8X5lwoAYKvHO6bjkOyYqUmPNe8XQD/ch3zJZBGMapa0CdiQ0Jur96Ts5TOYiNfz99eX7yYs0
lFgWXVcmQodUfTB6HEZU4rz4+Gzg5W4rZwULxsTcrYA8lAhHkPfNfUwJskLxSrYjaluW06FxDhVU
Ojc/Ml5gQxgpJUsrRJFV6+PIypB5Qln1t5R2IjM0YAgmm8iAHEaoqphUMCG2RQRvEJK0Y2y0EcG8
kNUWZajgVsdBeZ5i+gb2ADtD9aaLWP29xJBx4kz3WGI5Nxgsckr9kkB76nhdSNGwAbV/tpkXMinf
xDFhLrvqvDWMiDrvrH1XKAbHzxXde7rp6Wno9xom3hXzTz0TvU9bPTksGQ6FCMp0WUsJ89qfSbA0
j1WX0tdDVkTuNo7RJa+Oj7jRWpA2tjN6n4uVtlYjBiVswuAUewDMZQXUJDRAnh4AeU6XUQIfu1bC
MZxXmkLkNPCEjeWl8cyVp3ApAxrRBfOYqtVKROPsizpefCXbtGgwo4G92jEsgmW9tmnTHZ3nLVdW
Otg9RCAHurSRLKM+UvGeOySPyrKoOkgAVYQ5+V60ctjmjBjagZtclB2JERY6GxNvTuD3ZZTusqng
IihZoEjRkvd7hD4wvUsRQpFoR9c1f0AbgXHL1C1zORBpndT6TYK4OOUes5IAMC/q5CaBqfc0D3wG
Uqg6lHEktftMLevHYAvxzj/WOCtGR1iNi1N5EAT8PMoAJHjvCcjTioUyQcxHGI00u+GRYNgTSHGo
BbLqEyaObQm9PaQ//Tiq8meK723Hc2559W9ozik6QQVkYcLckuMBGod2yFrIBHWa0KnrcxHnSSWg
W7fm7hLoT3cDF/jibqUw1n/o/+AuAXZ96ld4sYvstdPf7eWdYdJcx/LkBBgkBqk0ZHLvTLWt+79M
/MPKni3MLLsTEQoYaXW0ybNoq2lpXbdTN+DmnwGPHC69yyo2jmnLcvA4ikVyOCPsxS67AT+82bUj
bwt6h5/gy8SxMCscL974FQqsrDqJatHIvspgaGo2C1VWGWDnjsBTV+lCrRKGFVNi2BEGSY0hJAwl
JayrJloMoG+ojXtKRAuKx8wlLizCMmq86fOVJOPL8Sps8po4ZXkAL+JEbJTfzZ6NukF58MS5jfle
Cp5O26qk7XE+lNUcysbKXGm3FzOFnSaQc2VSB1vKpXu+JAUKhxVX+9z/+8kdh5q0C+iXCViMW5uD
5pFyhGAvQ/7m5k5QG8ZIrpfaJS1e2huOAX1mfXhKRrYKFQphSPFB/i/owwll7D04bnA9pxC1rP17
LwFWhwpFyhKuAx+CbLKMEyGfW7wcUJXtVILnoJBdVq7RrLULQ+GX6fZN8s5VuzHa3LCBPSDwEk3X
hHfnZoVP/cIRQ8l1P5TWslcoGDBQZKWs8MWkRVHHjU/aaeFXyjcVY6B9bC+eHaNNE37svRG5PSsg
vuNFdNHdyIOIIfdv//y4s9zbIooXVTutTeW3vUKOlBhE6e+jSuo/7xVJO9ivnSohjo6UaxHeZI9P
njDd3Q1TGwgKpxb4FKR6rGVk4qkMouBGCzIbwZolFMCyTVf/Q4ykQmaYajWRgL80Zr3EuVcPdoPw
xmFnm5uTybGEk9Y0+DmXUJr03r956BmHUYzKNfsr859SxZYVE1jhhxhHL5mNJ6WYS+gAt4UldRHa
i1JN6DBDfKB7CWg4Y7yTUJHuPUSv7DV5B+owZ9xELwm/hfCsCJ/ol4vqdP3qm60aMFi9YuEkibew
NH0MO0PdSYycrtr+P5TOTVzA7tzIo6/bzEOIuQ+nho2YGDDJZAkdSKaPR9LulApJ7y8Yj4U1lSrI
zIz4H1rT/E980syYjU1OAP5NpvXus9HLkcJ2hpQFw/KI8ed49LQOFG/UCgOvvMTSeqjPHgJOhaNH
4/ZvOA4IpeytOE0Y9aE7r5F7783MMtyv0c9aAzpjq08G3cIa3yGOKUdqW+grvVI+wYoqkU+gYy/b
Ss1VC0OR06N2U0IV2y/0KzlXGuefLPjHuiHZTN3ZzohenDpIbdSLliX6geRRSBtyeTrw57p6Di52
Lv5zOAzPqfMtXBZeZ77cKkrYbOd+en6jSCmshZaQapaa6vossE+4ZXwXgoQjvKMhSzD/9aTvp42R
+ZtvcyjeJSySxC82krDCQGBS9ZvN3UG7r+qAu9ksSUaQkTXcc7KLRgeMtN8Sk8GPpWSBCfJCDTrm
VBpWpoV0CAd4abUgbKzUpFGt84jD1WEtph3k/1yomtXVV9WYVnW4F1cKGiVCEj9Jdx28VC/H7lgt
1yxcTdREcVaeyJ8fG0oilFNr8qtyDFdYLyD1PuxmITp607WE5aWb7LvmLZ444V242jENfzb+puNI
R6+VLw/QtJ6judxZrpyi8RiCWdm0x5CYaXLbo1UXrmk/QAHKlShTiQjMGALcWyE63wkFwaI7le8Q
O6k3pnwn8TRsVv47QEBVavB9Dgrk3B2CpjY7QCQh7rSsXwR/VKlDrfHO2PlBXEOByFP6vp5NXW7D
4k1szTvEQS6VW2zDj/yful1MvvGabjKlbq6kR/rMQLTp8oniZdCdBx//srFnDsvTF5nzNQwysMd6
n86cTe6jHgPsBrF6ANeFuhgjICpZTWHs/AsyUXsKMwMt7vrtdllJCXclDB39Wcc/hjLAma08uUSU
VzchnpNi9c524BVEamAUqvIh+ut6BRbJZRjH/KqqJCbv+LcKEbn6FbC1MT07+URoI8x7xEXEAWSj
USLBRivKE1SZQVjGWYD8K0iWTD8j3bStrvYvPT9jKp4rFFJV0jEAx3Jrg5wKYoQDpn4M2hYvrkME
1uaBb03s5cBdMyhZ6b+PVjT6Asz64lCTvEQksYRw3lGOtay+b+6EPMW8CytuTefifH1C14WVgZnh
rF803kBCy3qsnYzWNcntvE7Xh+mq6XLyNa7MKi4CNYYr9fW04nSKqO7xWJsevcVwzH+5ok7D8jw2
G3ixolvHs6KeIdN/naIPOIFqcnl17n94c3jWKOBOtHWCz1Uh+EQkSXquFq30SYY3CzLXAcChUkZS
TH0MjGq2qOgSZz1ke8BAuz3mmykg7JVgpzd3UUU9Dpvt5uC8k7PDCmgBuE9beYlBcOOoQV896aIO
HHmctbvb4X6xOY/Jh1WfoikAbhlIRHjujo637MhXA4UxFz3d8kCDaYZIWsSRF0wrXaymGzQ/xAbZ
0pbBudx2FSY/THXwmIbNwvUvSI2E0Xmfmtc1lDOpXhhGlUdVhBArVN7Mg278gBqyHqRNqyhQVSxR
8JQVyDiHShbYKEdxInSJubcWei0ECCDKNcRjS0gbbnwSqrgJ8iEr9k6tJ3m7gYQm/tOtnxAglFeo
gAg4360Z7XY6zk1HYEWOBS8sgO4TCDRzaAM0+SiI7jjDq1D0hz7+I4/1gwYBSvFtuao0rNpmk2aP
G8mqZLzFS0ZB+Ozy4d/YxmM5cKOFQLKXEb3Dqjfak5gEMElhyZzxHWWkRFRy09o3D30yvlGlgqwj
AF0kHJufMBVFK6L5TD/A8klIVpi1oUf3rscdGOy7raQ5h4aEvNwdWicSsOx1VgpKdY2DTsDqEksS
H4Z2zOMacWoxkQCzO+bXCyAMsCrE0oAgs5uhjV8UhI/mGRq39wiFoEiFdrsuR+uFftKMLzN+bqUS
edza54FAwDYTkCWv6ZPOz3i1UF5CBasAhsI2iIiUZnblvWVRhtKWFpuo9Mrp0sb7v8ARTtVME6YS
Qv42ryww1TnGrn7HRvhh+z7hdfmFCDE5T4eLYCJWLuVwsscNYSly5nlf/cqpgVCVeeevSQgw1gI1
paEFdVela7lOggRqp9HX5+iCZMZRHpyhCNrkriRqafCZWP62Qnmyw+rKK2WCWD8rkhTeC1o+OU8R
mpzNZ5fxJ3HSPlS/Ax1tTBAlTax7jOay/x2W3gauCKPlVq2eLsXL2gJwOVxp2vi4feOyLDVsjekn
M2MXCllaWIR1JqLbvZ2PdjiPR5pA0IDHroeIPIPPTCcBcIoFeHmyHe1DYQ3GUdUOFcvwC+xL/U16
5kpXH9P53ffPhLm0RD+9Ma00+eYNj+rm2R0KFcu0pavDPvrCthzZ2q3ZpK6APLsLax29fZq5hSvh
7dq/00S+x02NpsRwcAi8AjrZmWkMgu3vOF20K4Bx0jEs+3veMGkR0zAr1KEujONf7morPqrNoRmq
tcXicS+gbXiIVoVAHBg/oZ2tS2SnBS3I+IDflB2UgILyU5rsPZ1xgcYTWwQUqugyXyQffcsSYEGZ
FA/aqnE2aXh5IiTON1PKrUg38GEPMeTl4J9MgAXBChkq23XcvYn1F18s720bkxe82ir0OwsZEAWb
JW/XhP/j1g4ZaUemjpLWufewoaE0q4PApajKN5vxI874cMlHDfBIS64PEAX/2CSDh+63JRDeY6s0
+h+CyLB1q5GvlvHgmVXWaO+sJ7TDUQ6fbapuDO0hCwUA2jMepjL6up53BVXn0QkjLChj7lOBl2re
xNcJNCDWJgyWHdh02NiHH0ikIFvv2In4qaUglRw4DXCk1rfydEz8EoyA1cpAPZRhNm9SbwQpZOZF
l5XwnxW9xL58w9BjK7Gk98XrT/yIyVMkTdBQfTqAUD+D8A0bLPZ1Tdav3UGWV8Soq7LCy+FwJjVD
Gb6uJQsOsLT2TnFlCJVzdGTksZHguvJNXHlOjgLi86ZmCFsveGt8UAHxvvKr53oPRh8XpxWxzctq
WEIlRETInXcF0Rrg/xEZg3ZxWu/FDK+o/4+4zNupC5wJvYBAyEcIHltnjFyLxTWaTjMJIor5Ie9z
ISF4H/jzwfBqata0kErJhIyGog5hoSqyHh7229PJol6whVV/CPm5Sd61yod0HPw2Q1oMw0g/0zoK
JI9m8iI5PI8fjfHTKyLeekYE7RD8YZ7+P8n0XHW/nzY1kWGTEVhSsa/Q+1pV0E3xysDH6sMr0ope
sWapGElQIjAzCf9PHsC2IIzL+9vNvvzw2XneQ1w5PWNtyV9jYVoqIWXTUcI8cz3DuKQhBJPrlXO3
0FGxXVM78mPZZ+aEjeGKWEBNjO09YR2oOYki8MjdSi9tHX8Ek3mfZIR3ABcyo7+/Qd/2MYmZB7D3
upK3dHytfFqa4DG8vdO/2VN1Mht/OHmReuAPp6N2+LNEWrPtkER7w53zVwJ++CGFxfOx2SSJzUW6
s4rN/DGPH/3ZFTqRJ/ci053UL6q9HHOebd+IQKiNYc0ioeg20pIj82D+dkIUi8cykvCJlmswbTgb
XeM9Svfhg8K9f9P9jqKOT89EAchRWiszuQajRrXwB5u4qVcCJisegZy0hhi8K5JMDHiWxfUu6Pm1
EMjGPey+a2EaWvE4654LUYmt5zB0YnQSLH92qJiGxMgeQl/dggMSGW7YEP10LnOjn7zk2W3Y+gsy
SobUeFV7+q6IwUgAY6lvS87xPhLd9fUdKryvv6ZFPSfdpyrdQa9gb40yvcTshyTp/6cLV+PP4XwG
Kys60iEMu/WZsJXfdRvH1HavuPGojEQK09i3asrqS8iq/u3+kXfAU81u+6f8pqDbhsrNE9+H8M0/
Vi0y8yExnqDocX//zNIXCHAb1oBmAcnWLtdff6M37+t76X4r1f2Oq1oeXlJn2nKLRPyN/9zznOAT
kOY+iDXTbPLVUndT1+CLdJDSxNTajq+UqvnMtOnhC12jNbR3c5jHezegwn+SJCvRF6ZC9HUqpAPg
C0FGdEfSpFemQu7a5An9Y3CenxAC73f6Zf0tRR2lIJIRNPy9Sr52IMmTGoqceSAfcwPjYpzcZEdS
K92P0p+Ussbo9FyIzdnZoRIfBXBzR2dV5FyyRWqBl2rHqdmPE3x/HGB7TyTtVzL/4UDA+knlU3M1
4FcFMbCABBJIhOD6jX0DPPL8gX3CAtOQQ2qDKYgYHG8Eg1e+Oh507rPBGllrZbDKXizBSKwLy4WZ
0laZHjFZt9Wt+no/eBH3U8HoaAuxswASpaGKZH6Ouc3JANrYnQanmTea16c2Vl2fciU0UVt2Y1/T
ZjlZQFVktrCVmI73z0NuwQL//GxZWveZmTG+ZSxjptbPmua07/8PrwL3w/penkwcdefG5khB6xqm
nnWX3zwOV1O9UudW9NtHicMrJyx3vyUeBGY4v/+ZdDyN4aL4wSovBTTDUVI7HTygixlDO+8BpQIe
MP3vBrmfr3W5G6Rf9AmfXQSiEVQQh9K1DU6mEkQIk4ZC6k4++V4TZ4EJ4OfKrg+9n8B9M7jo6rdi
vdmQVTJdszPcAgSYufoOvxne+dZeL7zOUPIXP39Xf8zeo6zWJ/4lTXOy1/Du8KLG8wXu5d9ZfCuD
ry5GvPBg2S+Z0y3gK7FaSTg8KDVrp6ykT36Suqo0FLoB0j5h8VMi47ldECOhFWPoY4Cgtn5qe1pw
dfMiyBUFHRMeJRznDQFByKj4927WIJjXxrYZQbtkFxaU/GAJkcOVLW+Iq/klak4JhkbluO7hDVdN
MHYtPBN+YS3YhtB4z5RGLOYUGCuwShcqKXnM6tVFYyObgNPwN+9iy2N5HjdQaWh8sdk7JXVqSlXH
Itm+z/nGPX8YvbeHRNDtlguXtx1Dk6tJ+Rl+HACk3zOFXJvEpvjiI9VImjbebES0Ifgpw6iKz9pG
NhUIfnDGmsMuGPPExQqt0+x3wBo7M6K6xWreCCynAy4TdpsWvh4KPZUdvakIgfegG8Gl8tyM4yeE
9AvStXxK23ZCJmjIBjvfzJ7+Smhsae17U2zHrSvA3I5j6s/UfRcgBER61qsyo7jYpHp3qoqkYsGs
loaOwxkBRCy43pcIKrMfhNqhkxUpEkk1Lm1Qenbb/keqTmZOwdC52Yz1kbFl74+PjPFAYhy0RJNM
dFO9LDHS/P37yc5MMb89+k5MxPYso+y1MOxv9GE/RgZ0Q8MvYt+RhUxLczInIFoAVojY1cBLDbrk
JUyPfRUQaKnJ8uZ/TvFWyJhzCPiOxcLBcyJxm/jb0njDKeWBFOmZbSgkNHhRP+PdgsEfrqUw5QCw
vXm+MLc7kEFv7XIVuZ8voSmtkL9SxceQhJ2Y0H9AzeK5wWoOr1ReWQRr/SGXNjVb4JoP7bWJxGHG
vnD/jghfP9eyjLBEh7g/PNcCuRW+akVAvBfp2Z4hECvudM7RvVGklw+KKBj6YCwke8Gh3HlxT/8U
iiuwmRqW15i+5nwcO14zpi+QcdX+bFkohbNo9YzPR6dcBOhVDukZS9K1OxFREbIUJmrCyEJoohh9
kUK1qP9NSWQsB7vQQEnj+69H6xDipGD3dOFGbo1Nk13W+GqOjUk2hhT5xT45l+Cj82N5UsG6KQrG
V/agT2fhB3dSZyFyvrFqe1RLhryG8kxNCzpNe+Ca5aqgp8ef0iyX9N2ilwkY/NQFyxtMyExs2I+S
pi1SnjI/0UaD8zvuDSdalEm1Jn3Oc9mv38JDKD3WlDnW1qeKVjEGI1vniHgdtrH5uohiqm8+NqEZ
4+fpHKnQDhCAfpJpOhin0OCo44Ojb6/wA2JBqh1onRSz8p66KmAewU8/yy+3FWEXPzKaUvRndnEH
dA+6pQVE+8Ff1wyP5XjWTaOHjxnGypEYrmQ7E1xYhgDq4tOtFLRk4BgIbWxlqvTrET4kVWDpiKO6
k9lDUaRTZb3ECRHVtGMU1/NDaAgUlQH1fdDnGQTzcNW88U/Pqou5RVQ83h0TF6iIcIiq85RlN5Jy
B1bF71Ayr2UqQWJBBjQBIPMn6zrHswOKDI+45ROFhPjiKQpFrP1PuquCmwUA65URshcVrLgabMWW
NY7/ENFH6KAlC/Dp5e/GRBuIDAboBjOm+ZaSO4EoYAmutQOkmdiizyM4eWVM8Xa+m50hEigHStG8
4v/ww2sun+oUvPpeBR8A8dfIDPFLW8DG1nCZQwjdjFxJGISfnKyImLvDq+PsO/PHxU2QSSa8B6O6
SnlUoNYgGnOK7riGa9doKSFBDHMWAM9ep3Sh0yT1hjDcrSjrvELKKq+1T0ndw9pdBT6a5j4XdoAC
qijYX9kO5XujrrV1TiwypSn2L8EBDjXCYlq0qiTtcaQSkjhl1887Wga8hJ+hBA9+A8dw/6I7J7Wq
pgIEqynHFo7QPyT105rDPuXytfaGrntfjCtuzT3124lRc565JKi5AsEdM+afutvr2Lf8lS0CjAHK
Bot4s00V1ND3EdIOW3k1rC49bn2rsDNYKitNw/mC10N5+6RFJ/UnGiyx99uGpaoHuZxydWN8XZK3
V8UM+zAHLhlTnYKBxTPsS4OzElgQJ2jJBx13Zan1mbu5uwAsiYxQVBjWtvgZrEZ+8aj1nmYWh7yd
YopxTFXzIFVJWy9eeqP17UoH9+SclN7F0cd0Yoj0/VIeOJ95NwnRt7Jdvn7TaccQPGqahEjy8ag7
v/8hL2y/U1gk7SmjdVPj8JmreYLcR5gUTb626npblYXgVsNvjhKN1mbdZWFwhjBL8MpzTzZvckWV
gnVbLGPPWvKCF6baon6YMuJLHqknnKAmG2XBd8FH0W+WneLjT08/pFzA7+Dws1sQhgc6neJn6JJ/
pTq4bHqQdPw3wHQpYCx4PSnjWWkGBVd29gOZexw2xP7XzS+DxzqbjbKt1jiRCiPahrMgUgxCvjHi
1eYSLRMxDKLwkInMv6vQwHqY6K/Yilf3ZvGzJw4LZyhtdQ5PVB8idDeh63o8djNpNT+whHmqjKpZ
SEO80L/9b4oGn+5tStgXg9QHSsm9nDrEcycMdx2UaPyD4eFLwnGeodYWem2Rtri/9Qdjshckgyyp
0OVl2+OFhOV0D9BeU1QLnK83M0X5cFWRyHbhrPMAXv1WQXA8LngQSulpLkdoyAYxBy9CTSQEEtIR
yZi4nrRZATIGEXfOI5ysW+0JlhZb5IptOmX7KyH9a/ZCX7lN8GmeEH2aJtNYxH7eyY6QDP2bP9Fe
2XJPTLrc++GBnLUXAqO8OAJQQwrpKZklmITUQKQLl86n7RCNV0m/GfgD7LRirODjIpwTFJgb6Ibw
y7J1heqhlsoUeUW0Yv3Je641akqkIpj83q6CsuQsM+l43wbFdnYBO3GDlwDzQZB23MfRqYRxjWA5
3q7Yode+fkO9Y7lZs36TZES9Uhf1pSqyj0HCg5otHDhOmVguMFlw+FhNVORz7oGHLb4w2snqzw77
UPwv8XjPxqBCYO+cZTUnWiZsnYzhlDLRXHIK3NwWM4hlDrjvxK1IiAjQ45bMR/8E5POxG1J2iXjH
uXX+WlGsEsonStovGXz8yqZCb0fE1x4FAkaqU+1+xhSuxZcUx6DSlqV7DU8MW45dFopaipMMdx/J
3wxiVecBjctYjFXQlOkbBG6tt9KPZiyLXS5IcKvSJZy4CUTxX+XBWbO0HJ60rXgGa2nKP8El/z16
JrTsJBc4k4cKMjRswUH9Tmp+lANQ/Uu+Jduk75RM5uK4zchyGmiKJSr3ool6CIfGz77F9QpVkXam
X/Lmg2OjVVdZ9QDAPCX9zGleg2OWJZhDJbRHivOC5UTXTzQjl5b8jbLkuj4q8KpIYNe9yauhuh0k
kNzYRvVbfG/a+aIgsP1STFEcOtrXN/2VIrjataX2BdIt249GQvD1SCI2whBVX1cl0cn3IA34g8Tf
oPz7H5KgiewhTwFPverpH84wI+Ze3E5kcTI1+UA8IYRup5WGCmUmXwAtzyL2NruoR1fWgAFKi9nT
SnUYBNyuaw5toScG7InYiy8Azpbg3D90IbeTndPIs5+edZ/pfYBuCO47Qds4/b5M1epRiySgEYHb
DkSoVykFCC8y9W1jfiv91fnDLw0zeROxvvY9ELCV3jtW8dPkW4T85HZcjDr/CUQ8fyfwQR/LPTlw
e71TdGm+0HJvpyyFAOmgiqnUm7WYWFt4toOSFcxNVoUq66C9qwuEDDCbclOJsMAF/Av+k1pMuO6X
OXiWb9HM1mxchsNpmhUm4srmoln+CUjznY2lCyLojqKOonCqN2i8/iS9E/JkLePl6K5D1Bpy/o1W
kpbL1e6QHxSUfJM+HyujOlZZqutAXNvE0Coibc8BSMWMv4OAcPVqE0+ipquRAyHq1E30InDswclU
W8Lo1nVoXkf2PkKYw8F/RO8PT6RHq7KEJIcrJRyjMeiQP4NCKjVj6a30pR7ZqF1l2SEpsC6hhdPv
7dsc4spnzEKScAh1gukBCnxlTX/HbrMH6CJjlan1pIJwFa8OoqoRHpv89Ios690CH5A9rBEcyVTV
TMQF3KwbZsKzR61zheUpKxTUa5rtTmPOPHe7pmlAaACdGHNzyfTufxiEnhVt+RddgqSAfSfIzJZ4
5Xaad439z6CgtcECXYagt/3zhcl3uY4+RULVQCIQW/eMiLVBfnUFck/n48Yr5Yibph6D+5oV1jvn
wBuHyMX+3A4aYZHuW6JvbsZRG5nkpYx7mAeHA4qkqoeHV3ZCTMPonWu2qYUw8xOueK4zyba5V695
qEQ4MgTiiX3caOYZYRMQcqB43Hb7mb2lKahB9OQ/cpfDaBsmxyXUKft+9Iroz0ix11DSxtiWGwNn
keJFl7/tivXAP/oZfArSzbyy6o92ErhXEaKPk5EBKx7d/fwfY7Yq8FbIezqjJJLav/coY5XMxTf2
G/r+4a+jsb0M2DBxSQhiDaga8d7IiIDYsktXdI0Pi/8F2Sa1sQGeSp4HNDrAqYPbdSo1wBLhUzpg
YPkcr55x4CPQUpXYCMAJaT7Hv+pTtaPLPqx96size45lPQTAxWynfHRqoNtbs4lADGPKQM9Xn23Y
M3P3Cft4VSXjdGZL4FzqQaxlWiPIiAyY7QMKWDL2tbaayNlTF1zNYvT16SB6CD8hxTixH9TLqDbc
N995mvkOtxnZNX16ToHqI9OyD3z3nA7A3gTq/GO834SKIDcEmNpa4TS/CJqIgALt5z4us3juia0y
cgcWF8dENp/0MdPnxoUNGldajNmCwAkSCbcByiSRsVR/QQ/6NcMM+euovm4ZZdnGM/6qMFm58VhV
1jA3XJhmqpIkzYoMNFuwZiWXNArGZZMR1rDD99KgMZE/+XOdhGH3V7y3fG+oD1oaq77Ivt5YncL4
1pGHeLJQCG85LJctaeTFHzNynoNhgNBtD8t9lQTAs9v3GaVlCGS0osTt3WTjgPLQP5SjTNfTUpHa
1M2oGCO81+aZfLZPWbkSbN9g2wBgqBfVf8iXeYE4RAJp9KQv5Qptq3tk3bclmFA1zw1DRAF9LHk6
nV5SqzV+qNp93zD4jRtQQ60/UY0nbS5SMZm5JxeVIcmPVl7xhZ/6u9QgtTX3Qpa6Q3RH8+zqCJW3
a3OMpMyB9744FLVgT1jeUUN1b4gQbdpUSa1n4J+/5irYHKEZ2REdSYHY0WS+d2r5LE0U4w9AV7J4
DcpUbgS6vRgeESVpkUCP6kjkBBQNAjuqv6NEz4PaIeOnSPB8zluTUbIZWfsvN+nMgxgefH3PJPjZ
w1qFE2ko7qJIxyXTCwrZ9Mi6ED1+ZGBSk+fkUyx2AB6CBAZnSGgEOH4px45QMgo96G1Kv+otNbtg
w0yZHbRLhm0VrsniUjxbidj58anWh1IhWsI3JrNfM2IY1BFokIRq6YxVgon1J22AoQBUoYzYow2S
bdRLBNvnrDhv/JT4lNg5t87PmmYrz2cqAB3w7gfNv+PC23BgvMmLT5zMTq7yT5etUV+3K8AV06Eh
6OT2Z+vPoWGOhKA+uz5PqFxDPHN2/xL77qI1tXXXR4vu0AI/EuLlHtwSUaPMi9EsTBL9orxvn5q9
7tjYQ52J0znddFuF1mlT/l+10fqsn4JCcOyoYq83JPkzHe1HC9nGeYZoDRoptHuBHqt1Iq+mYw71
3q+KjYVFNvNJFNAEcwTGIpLdRYRptNUtoZmz6aVHN02KuL6fHsIdUeYI9EdclBntLl+QpssuVAwC
GAtRYnkV/lrVCRdLM2wgul7KOz0pkGfGh/wPC324ySJ5VSxDt0zdJd3Omp3unPZMFrI0p8WCKhvD
KVkEBBwuiGvmw36/6D5TFBhMFR2ZW27o6PUdEBx21wxDhzgotZ+jk8iK3K7WBpTsY+sChaMcpYCy
79SeJ7Gg3/ezFCgmcFulykKdWvE+lQfWfdK9QMSWXAl6zuvxHiRwYMOjiWZhAAPUJYnCY8OwS9qB
LuBMCyjQDf6WGwkoNhzvNy4hZQtz4Ria8y6WQkic2TiZyquOwDILyhdeJjqT6b3IMbyqzdCMDGwv
+bsEwkM+88RRSOltaza2kPYT01JiIMWMFgTmFWCMdbGd5W7gQRTwLVDP6e1B6L+12EkQ053IApQA
cEuUG5QTvWqz1vxg4VQBilC6coNvr+szU/YkBiN5C/tHUVkrlHzF5PaPA3Q5OYZp7OaPHVSZuoqZ
u6tCIerFgZ530HGkyOUiQADG3L8XLYLWHeWa52uXhmbPXFeffIyrl/Zt5BiREw/SftvZFKpKcjXH
4OPb/PFehlfE4s0lemVWaArypZqXqO9yuGutsKiT0Cty7TCpjh1Bvt5PBMT3Wt1DGhOGtr4ZiPqo
23VA3iCc6u+6QAAOS5pYqoVNBtE6KDPBuqSCbjCr+oAlvhhUXRWv2JDQZRSthDcJHR5XcmyPqyWX
KqeMSLVT+y12Ylonw9aenv74/wUy/QnkMSvrLSsprbU8uTpdLO3hRNQha+2xHlthvlATn0LNDx+9
bibTrLXtdrv3mC0zT0y4fH8wn1xmAuycf9yLHstn44UvEDxU7GFK2JyU1DpAV2znABAcJNjkqCpe
OW9ISvEaIZlHWc872GyTjVrPkZMgTALG7ctsCAeaNuenK7/0TNVyG0a66wSDBaK22H/suwHITiZ7
XktQsfgFdFB/IW5gz1x80ERrQagHK1HrAV2TNUv0cC6+BMZl3TZMWR0mp0GumXuJ7oNDJiMB59Up
x5FqYIL5C9TUWSm6N81UoEzaKrrUKTruE1FZkwKFc3VqTwuI7yIbgAlYJat9E1uGAMmQzSkf+b9k
ruPhWkaIEAfu0KCOFhy2HSaEGOXhy+SQxy9a+8S4shyLznUxRWNvxxd0WZ8Y0/uUaAA8HQLFu2mf
8Jba57ZQ+cv3moFZQvZKp5Cte810oYu0VujFzWZ9Nx7gzDf6l+zofloY8VnF1jmXzFg45PNnppav
Pm9Qd2WbVBWBN51WCaSyhF39P6a20vdtNDKPwEPRyXz4DIXWmE63O9cwh6svXu7dLrIzFFzAmGjy
bCXLSwmIv6Wrhe+YtFS5r8ndKasDzE2qly7K9MIf4LBgI3bL2/8wLmhkxtj+YjzBxjHV2JX0knKz
6QE/VAPLUHlSmbSHvBDWn0YqoK0WmbvoI+LClJmz2Yn/RS1zbgorTmBOaKUwd03/gNbyKSknP6Du
gMH4GQTupId71qNjC1yengWsE5BLHEVEJejB2D4uQxv15v5+BeCR4LLH1ZYMZwbEb7svJKO7yyt7
yDfgz9oU8Ny2t7XsJJVAQBj++2DM3N1+0ZF6bdRNTzVrgweopiLaYxxifUfO38UuO342ZSRJuKiZ
D8z5J/r7dFE5Xxoo8DOVeCflHcyiK+MITm7muHC5AzdKx4PkwHdujwDnMOgryQqz2MhIURgxM5Tj
7vHLf9iUbkZjvyic4/fIifNZGfjSJWITevhwSx4Ny5qdnj3E9LAWDtTtGEqYUchbnfhnMcSmuA4o
4Tm3dMWj5XA2Boj2qcbYQDIkLHavoTiZuCeNZu5i524NebKdSERugZt6X4mt6xuWFtkyxu6bA+xP
qgrypC9TfyGZDBfQlfEO/eRkIrqmLR4C5lmMd8pdefk2vFnojjjsONqTAZ4jRYXwyvm2AKlOkGFe
WeFMASq5cnlh54EoPwiBiUjxLRnU5veD1zDd7H28ngmzcRnHIfQfHvN7N47GxOOc7Ud2xjt8bv9W
+JM2BSpZwD7Uzh/f3nh7H0RW2miHuPTiRyqBWAimOJugSWww3qoFraVv32tbwjDm3lODJ6OzzBY2
KAi82V89JE9St7KWx9ke8J3z1qi8tcBHk79LpbfWR121rOqytwj3K8/xeutNLybUlBmW/xbLnI3n
uTmFiCdcOS0aVzfFYZ5ClFuyFtV89hDWspiNXoDo1JcSid0BO3cEOai2L91AhiVNrIOiZnd0u1RI
Z7eBPBZqmAAhntchklRNqop3zrGTghcyMpxMhLKeE3IRdIAc/DedXYAf7CvsW9akDjzLtIbFBFoP
bUMsXlOVkpqQiEl3CN9ETp+nTFQR5HYVz2co97OWmslsfmpQ07UfMkEx7BVeVGb/sZh42EyQ5/97
SLY60oG7qYRLZWr8tr1FGrQCFaXefeH24iKaR54hO6lJkQGwUXMKYBbRJHKzF2ePfbaJ9HSe7tJE
k+xGV3ddRcEFbfzF4n619tcSKjCakvCoPbeN3Y83fmsnnAntVxp6AJtAWzPt2NecVsi7RGFSwxBS
d32saA7e6iVZP5VmdcfdChshxnufIBbNZcc18Ebh5SSwnmV6cCSltQ045r5hmNNf0UCILRZvgc3z
A4dfKXJHzncR3iRWcFFZwjax/5VG7i5rOJmIH53Ve9llpQ4pcK9duErDRBLt/hX87Z4laDmMwypP
h7qyApfTWqDbAUWB1gnYdNhk7c7WYeUzsa2ANSSwjmUSttjoDGzW+BlwrRThu4yuzGtG2Gh+CkqQ
tVqowHrF9ZSc8MjGmo5eA1V5BKBs6vJCNb0yFexwI0Gt54zIRBmWfkAqD+RvZ2BQiop6JjoUHmEH
5G5zEgD7R+NXEyf/0iABx1qBl6VpclZ2tMHYxu+zyWUAJ8G0hHyBwZDHVtQlVGfYoheXMOKhv2+3
Jv0mgaDj03RgKExrQPkWAlREquyARBzgIOzkdRUWvS3TgsUQsmPMPKREwaOuyisbvYMnBAllJVLV
4I0+7u4SUETVTJHu4k02wImr0Jt2fjNsrvFSyfI4fbjKcgJ56Wt+3+36wmIg89mVnwY7oeiHts5Q
xuP+7/p5GLRppfFtlX0MSPr7W0PxwlcbVKq+WMPzdWgLjk1PNbi4lm0d7PM6Ppt48/K84LJ3Z6Wp
lKgkQNE6aCPVUiwZ/tcXHMFs1hiJuQK38q46fZCMCXtLuSfw/lYzdz/nWWfyC/+WEaFviIH0hBCB
bg9Mi81UU7wWU4lifDVpEI+WPenxA38SU2eBXgvolKxXLJQhS+gbWei4lAwkLdezoTibzHsHLW7E
EEP5VNIVyZf7j16Og+EWAzN/+XiOTHvYK7K0UkG5Y1ElrV2oT4l57kRsr0auwFJgvphYwSirsoPD
nX+JzZ+5h+RJ8+M/dZgFFb9CdnbvzN4xXJsoZlUdjsAJtz9hVc9oKR+WGD+ZsZwMFnVzn5G3F7x+
KfcQc1cO8NZJb5GljoJhdAEJVtgCpQOKUcAZ9frDrZe2e6jtbPRHe5V+q6Vc3CwMyFETMuQprcnS
EMzsR7WofT3eOcDfjnXh8i2hxkN9TekLtv/r+CbsEnZ67a9vvL8M03APSFqv5UBL00ODgGubRVkt
4aYmyHj4SDS8KDFavmDcMJuj6l8gLHmzcVjwtM1Zy4ufpzwoJPAFCvof1smPxdAZYEefZcPJZSBb
4sIwwHcX3KrySfUaSd4Jh8ri8oJk+odwb5bT1K7KWp5nyIrCKCV7/Z0pIeatsBNNz+NDjdkEwp6j
YdXp0hKww528OzBAM2LeU+2CuQNX/lIkXWWDBTB/+L1bBNWzHADawTBcNH5MmGP7YOz3qVK546qV
D2jkgRhdS4Q8alttakkol8DriLon8Mb5p2yb46WsRdAlDyBDcoVFYk1t72+v+2zN4IjCsKeuqVoJ
RcKukP9JGIqWygdxTsrJuFn8ODTwT/5Y7Li3KFLYSvHujlksd/WPsUqMd8PaLjzMIR/f6VehCT5y
iOp+4iS9ncn+BbzW465eIri2rzoWYYorFqA85qv1O40iNOYp7o1oM+ovvTafkFdjlixLpq8NULEP
uwsswS8bL33QpSRNodfTBrqiGux6vcU/W5N0oaHwAeGplpJ/8wwTv3V9zHrmJHuMINB8Cdez72D5
BNYkdiNQYNLfRVe47uRFnIKDpv9HKbmszEoOwVMRqF85GIf9kzcdsXz4ATlgZJiOFzhTmDxROYnV
FBPbjOf9ceDhdTzrtGwQScN1dCeDYWPTka5RJH0GKbvPQGQJz9uG7xJzuaZhMmxL11kFFVyJGeLO
h9DxGxh9vktRkmuUA65bEyBtiHyUZcO66Zgw2MUA7v61ZBTjpDdQT1XKM9xeTt+XZH8GNaT9TcRa
5NxdqJXUkBu2I6/Whqs/5m8Eg0CQ4GS1bewfhNoPCMG57udK6ggwQe00RH+MGoVHvXqlakMHayhO
jd8TN0IcULDiNzmkm5OkH+jUpH0hqtA/8YQwaoCCUu/YAYpj8viqlJiLxUYEomRL/4D783Ye5lPg
dHaex5+9pkzDRespXV4u7LvujwKn3m8TNheHaC1eM5LV64HRPhFzkeBGCoffXDbFIHCEPZo+HR6+
RPbJ5pzF7PCMikWZzVkfNENhaCCBWwDEpYXlYmIWFEmDQXBgW94NnalIXMZJPgDCP7NSGsyXLD0q
155yMMrXF7WJic7ak0m7aFbILrj9uFT2pnEVRIFC7QA2l9OqaFM+vxfbyOWYK2NBhnBuLuR6kKoA
CV5SeIZqlqwL3H+sbvpp7aw6wXuyxDg2BSSEL7UZPwRypXpftH4XjuvLxU/YazrmrW4BWm6B9ByI
iDjM1abgjuqe4cImrrB5JJ58oN7MhSOEY+Hp9a3+CZ6S4mx7IIHwPmVx2rrh9eP+w6sT7KYP/bSS
CmKzLq0ZawRH6J1nyNPg5xj7QfMPFyHtr9ziHdW5YMZuBwaYsiFdP3V69nXpDSun+mUc1Rzl4Jc3
CPJLwpg0kE6TN94xeun8AILqUE/LLsAWxxC5e/lKhHbW15z0bdpBpum43Kda/H0VZnQujWYB/UAa
uMjWU/fnzke2b1fNM3O1K7giRysXJ7rAqif/TLfFhmMa3oWR5OqWgieJqpH7vCytjIKR9/xXMs68
/oWCtSsxb274PZMxnYd9QTKMdBOTHd0Ii08Yr1EKbyVQxYp5LaNZMfX1wrkIzQlG/SMUBBxmH/vV
tlu3IVv2ezON/eEBd+3Ygnt2e++b+4L/1uDiGqGsm6EOxlJOnRLFLOMtSr0djAn2hlbUCPKK7RLD
g42uxEc34Wfsu4DOsGhkGhNuRaSiaXF+OhlFQnP1q3hwHomN0cUmi4IEG9J22ECdOKAWSBujmPEU
P1rP4wRVNWWbouHS0tu2+Ojt7d3asSOOcRMYjG35r9ini9JE4y0y7+75oyoxdu6UdZhP2P5eNe/Z
wAiQyuG7NDRyA2kTh2QRXWHjdlIqCo9L1gpDrTCYvOd2cEHWxvWJgwA/mYnlbwDos0HTyt1RzxNR
5hY0JDrrx6StvC0PtcXS+nhF6IbAazy2XTD3ESDJWb59eOm2D7u4CPk235PQofli53B2f4ljb8pu
uCQpF8S3TPTWjVe4bVPKWuAmJcgk4tvyfO5FZ+lBp9772Hc7SXHrePMFOhZ5gFU1buaqdp6e85Yu
AQ4jtAEFqZj9LfdS/gmKw7vXlQIDHOt8uJ1NuIE3UQMH8Ws8XtMGYBSFxGraFInR8gZPx3l4v5WV
vBzRIwmOzafAkrm55wuiAY16iB3q4xvK4Hshi0/TXKjstBcM797dxxoMJU3acQ3NMUYOD1iid/3p
XG4ZltdAwfLUGG5lhuWdrY6K68dheUZwMZoLBH7l2udTuZA2MiPyM3FRdJBwUEJ+dIPB3yDm3P2V
gAnlV9Jjp8cSewlP/FFxG95HxmTFHjEFGFHky7AKZL5bLzZoLEzSUhEtoGVKY58D2xBeKDr1DTku
gERMX8MM0Zmy6x51hB6On72RH1qbbXsIHXHcE1eo+HU0Hg5XtM9XynuGOeLPwPVOgyw4lqMunVlw
DsHny9w0iWJp76WFcTxlAp6s2JTaKnqDzTO6pgBxutK+NXgdPCJFHj5v1EUDpTIXrUkG7whIDXD4
D1qlcWMD+/NdDVJBdadxQQNW+UJqumdt9TcAu3zSbOr3v0I3sBnlK3MmNfumNQZHlXkJ+JAFxf37
iTHSeRv8kvANVuETydata5CSUAZ0dfQ8/AWsYfKA82ystiXBNtqrMrouAlKsea8JxEUva/LZosLc
stFKeiwf1esX6yF17CQz9fAQsczhoA+cwt04ki9nOC61YQEmdtqMC3Zt5oqH1WMGlzrv74SDqS8+
T8V5/s0/Pvxg2AfSBQOMFEBaww9FNRD0uhnWzEzl4a7hdPhxDWN/QnErf5EVoivgcXylTnOqC8DK
XkzQ1pFWwfQbC+WbQOifh8tafLO97IZjFauF9hjBFuR/1h3CCw76asgQJ6lYWZI9KEdSryQxN+39
XYd0EPpZoIi3Fhp042WTZPgg5RkQp169gZFDisjtMrtTfKfWW5HKacpzGxCX7y/Kzn7NmFMU3RyY
07ZfbgpQ+Gv6ZY0AC4QTRczVDjm05xCghFzlcS7aB4t27CaSIlREekNfrGkfFANVAhrzVj+l0Kaa
4cZrFKiVvJzOFNqLg8bIQPYy5tsyJ/kv17Kp9BMwOsIihMFZmBt1ap1ljxNWF0p3gYJFb7mw8v9H
gdiiQOckVbN7UqgswoftGfp8wIt+AnouGqCnNvbwU0TM8yWAKqRQqd93PYZrAXG25kFI5Ia76fNc
0boEGW87Z9+X296hR06JsJW5yF2NoX9idEBnAKMQk0XgR1f9bxKt7CRCrK+RUfZi/GlPbDTCvZ8M
2/TeNiJQpSdK2e8i/bzgihyj2thlr0DxNw8GkMOxPZKwg7YjjTjPirgUe83TwkrFcn+nMgCj7HVp
3ay2G/1CXrhx1FSxW2AgJ0lr+QjSNKi5SHbD7bTVEAWWg1rvGRXKfW0eO0YoyDiCuwWk9Ow6NYh+
jnS5EvyS7lItce/qtzXzw2EZw04TM66avTSBzhmHv16cH+uii2AA3OUFTiJaXChymSirqNfRjg1e
o9T/c32gqfuKC5ZEBsYhUjJxW4cKhvrTvGjUh7144qZ5LcP+ntsYub6Y7z9Bx+utuutxyqGebzHo
iIm2MTvin/mBnE7mfPy1JYW/sLzi1ehV4LIczmEeOFNsvvz9koevDFLHKbb5BlDCARiAdO/LvvKT
ym+uHpusb4Igrz697cMVaBWQPci13uZsbQc3ROsbH04G1sallkREz/uNWhSGe9UEm1QIHZbU8x3j
TR81bgdobKVJwn/0bj5j+TXM9Sel+IPjnMdcyylRZu18KGizBCVeFzC/s9msHnGM8R0lnPvYD3Z5
xAM33x5H3tBEfgBJkIGXRXtvFFgY6q3tdMtsEhfzU+iF3ykXmyn1G9uMeqXaXChq/Z0MeXCLvjvD
Ags7g2IrS+AbEJAVdOxsEMzsCsvysdb2LlzH6n49zcMvR3Rd34+ubPI8X09EYHcP/qw5tlB80lfg
Y/XExZwHnu3mZKeS0NE9h/am+MbMxkaI2mO0+NzSR97FDZUBK5kYCF72gJBKskl5E0Q4DN1GFTjL
cAjkFFwdLLIAX0NdVEh+6c1fJ+7Y92F6VaFsyCGoiofjOS/6cIj8fsu60SZUhXxXXqLTBPeY6B09
zf7GiYDrhvuJlG9cTeb4d1bAaUzUjzM5W7Cr+dSsUWNn4+m9Uax9Rj3vZwVbGFhXe8yKhCn3HAtn
0rVybWvufOoqi/9Gzt8R0c0cq+4yQ/MYRqRiY8tKRxaTcf7UwTz9hKfS8wKKvZaQxm/NzesK9C38
+YO7TEA7APud/qlU5RP0hJU48x2CQxFMZcC4eYloF5RNOTEmOqv6+L95Ekr2RkPvwK6R9BQ/wTcF
2P0/hNVNWiVa+g8qi35dmq7G4TAObkSx1e6iqEnsjdJ3IcWIpT8LhUAsR1dJRkgzUOkoNCcP9SJp
IacUA6D3uR/x6QHudedQ/6l9tQViju1oNPE4bL3bMnMbunD77NY7TjAHOJK3PoKwMxIiJJrNMutj
BjTMNtur/WminHFWLa5WLB7piXxdfCHBv8uc8k6V2LsfvC7oBbCEbek0WWR1G004Lof4jgxFPAQR
knIo4Xh5wIhkdW2wCHyoo5WtUHhkH9oS8zT+gS2DKoK+l87bGIW44G6w1+TgnMjkVSn778b3ic/x
jRWSFHZs1wydyyB/kA8V1Oa/Z/8XoV2vpeaO5ANGYzMoZF4Q3AIMpThRBqtGmi0D9+UhIvfnoGPi
langiUFv7E6UC6rEaZM9w+K1zBAl3oM4rUaRn7Ozryuyh+kyz4YZVg/thgmdQXPWgV4HisLFC67J
xdl2rRWxh2NMoqhXlN87I7t+L0OdNUDBXxGexgZWY71IxYdSGANV1QvlruWSJB8VCir+Ov1xRf42
lvZBD3y6nT/22UiTKoqRhMMmVqEBZpWPlctJzbmYTEv1ISvd4m/GKAL7pMF+oQ6lzLKN+IB2SDqQ
fw7GsSwVsIL5r31/mAS4gkCax7OOcviKnFD0/WU6eUk/XmtSFPutX4Stz2BLNx+s6noTI1yZQomd
HQSDNJzW3jpCwH4ewEvuMNrGwWuaB5IsA/lJxbGwvcgtRxhOIS7IM3/X7PMoJ9DyfHsnB+mv17xf
DrSAwFFIRTtQMQdkCAhpifs6p7Xb5DJ05pe3PfZyYNqkRmUWS6Ix8tKRXJ/E8c8O5Wtt/qsJRLBY
SHAsdiYI09UYHorBwnqyaMbsVS2T/rSt8A4kHHCWvb2xXNN6Ya/koxpe1udjsnKtCXiGAHgCKvjo
GpXyjB9n7weXhel0m6TAtMKuNO1TDBs6Z7sDj6eRiad7vDQSl+woazfTwKsKCuJRG1Zlm4BNRW49
otXoWY2ciVgBTqC1O5otST3kZ3wNnCbUx8kvuJxP2CEW+rrXJ5ZAqkIA8WYkuOHnBqoTOVEY0j0P
uFpXakBO2gy802onmoN4XU0Lx94MEUFbt/T9jOZFgy+H0Hfw0c4ndp2qKUYfHyTq0T7iEhVVR3GH
6zFRu3T8NTo8L7ZUX2c2Y9eVJoiFm48snUMRFujDnblKzIyl/WtpeyeeRxJDrJenLcUb2v5/kfwT
UbZzxUeXP5KSewmd6+/OBT6LazqLQjAXtGGAsBTooxyH2RsTrwxdFNh3n7NIMIdPjOgoKZGCP2jU
Q0jCoM1Ls4lCKSXJu711mLou5rRgdNren1oObVIxNfhnaT3coexQTXsGhfm5emtt4pKFct1LPsQ3
zUmqxOkltRkIJyNGiLtEq1QzNpltCe+MgR7VtbOJZQxYn9BxpY2jOpOFLsLlC9lf/WGdj0mpEExz
iAD+p5KHUeCQMSBaJEJnD4gCk+H/GMTJEh2DpJPSRqQpu13Hd5Tbj6Q+0S47F6okCWs8qvkK1Vzf
L08SiYEOWH8LjZJyw91w80PY0aXxhpNMIUmPgrgjly3qd2aGQCbJ/z8kcmQQwa/pNXu4Ai/lk9Ug
0XZDvn3rfLhf9Dtlpiib7F33pIz2ZgsokDj3Kufqlvu5fdGE6tRx/JxNbx9vGhfdihm1codwxq8L
iP97nbVONUc8F9msKoQop2qr1L7K40NqtHX0vUFfAmEDHv0RMCsIC8UIz/QtKnCxteqAi6fsyMyI
Sx7AjS3nSUZ7CLdDxf1Y7QL58pkNS3IvC0sGddsL1qtbF9Uf9hoslJP+6UoiapBHvU3egm7mYWbP
xllL5P0cq5+FnXeQ6uYFigVsbiwSrUIv76OH9qcJrUvBHBTKPqiYeeCrUv7oEwfUhl+YHqlaL39h
WoNZf3okEeoT+R26BZOmUgeqIGWH0QreiozUUtrSsr1FlekEu6RuQDGAT9q4e+GpmiGTAVrJVrW2
nb5222RJEdt9xorhku3fYXlnqZxQ+hvWod3oiedHgIWp/FqAi+nuT15TOSS54BW9J4M3JwpsahAg
Ln7WUpuO5jiuRJLsTGrkW2YPD3bGgUHfaYL/q+ap6qH9aTeiBOVV1XE9/T3A41RCSjO1wFKFsnET
T1E0TT1So6YDQt/RpyUj1g0yDzC/W9fPEObYrOp7NMHrGS85vJBRtmaeQ+L/ROzh5PVdO/2ulK4y
HBLVwMqZ13/SYVECLxBYJRn2s3lu6nJsU0R+AahXah8eWW92tyzbZhp/mfJsLyqkEUJDzxKGhwAe
UtRjgdIdlVlqIS7OBX5lDRDROUOAU0hJiSKvXcAEhjRcP+65mjK253v/n5qyqYoEGvbbjciFvgdH
hhjfaM+9rwibWOKhaHAL2zICl6FGcJGVZlURSBillDwkLvoYu/TjkpHHNDtpyIyEu32czh1bKgzI
ATSVdF4J+s9BA6czgkWSnL7zhmXtUTguilUZuuFPE3tQ3y7QwN1OscE7BzXsL07QnYVdgnj2zJfg
W7sAp5dk4wJ06meyWQv0PUsdzVODlVtvxi8o3kIq789x/6dJubDGe3RJepSGqrPNLh3eFiMoZLrS
3629MQ0x50l0tblQrizEAX7zU1QaLuzJzahVDvwDOlFOMxuwxJ4mS/tAstbnbouyyNDwgpDOwBUL
tWDrFO0WiRqL8BjmaudBoanEUWv4we/C/ouv7ZNO5n7BRu5C28E/Pr9sfd8S9dOzw6+aqxgrIRiE
iNBiDfM247YPisQ5yU89nxokC6lZX1GhP/jijJ9A+dwpWSTCQLyBCcwY4VQSfBJRwwa3t13H+1OS
MFco3aR7Y2A6CpbQ/8+MG1Q6Qrd7oX2g2lGogvCL8TydK/9P3Ce+x8garEgBsJdTgH1BnYha6XvU
2Ewb+HGrqt8852weJZ34U93CYT3+DDyr6FYFicDlelaocvv5BMqAAqD3P2D2LpZBkbm9Jj3WBKKj
CTp2Ixo6AEIyDGqbR16QKomUYZDcIN/vDpWq+8BrGMXk2eCi540GHMXMmX6J7qm76L7HI/cTXBsy
LqIDxn+Fc9zP08dOcq903UdChOrJnokhF2qx84HACdjaK2WZwbfErz7L3226v8O3ybZVqEFg5/av
qL7ujlVZK4NxCtplwfL8VS3n2WMlvUhcwJhH9/qqQabE4T+Z3DNFcpMkw9znx92Iyofa6PRXa04v
BQo8/kQLvmLGKuy3MujErFKjGWlgBgJLFl4AgUSD7BlNOmY9aFAIsOmXgsc+JEoT91abhGLOQJJh
91RPuJ5IWd6BS+5FNtN6+WlEMKFDLGJ+ANN+t9FPrRq7IDJ9z0eaB/5IKLIW/BEkA1WpCYK9tgw4
B3Tgt4d3tVVtgO5YVirmLMuyG3zqbwTZLF8bjru68ANecuXhtgWwcgMXPg6xRtxo6tPe8Xc6M0N9
JyKPcJu0EIQ+ztSJwKsZa6FzmW/YdkM8hJiuHoGpAGk1AK1oC4cF0EhuSt11Slnd9ZCeOx+ytI8Z
GzZ62GMmBYNx8d5gNzDr5LwcKGdVVVDA3/6iRGd2EOs+yrMeEagFn4zm7yKIo00u+SXjA412JsVH
IMG281V0etVT+2+XjEur4XkBdMscASuA2HONG+L9o7UdKWUw3aZLAA7Sn/Zs5NJFVtOjg5oY/Ony
yov/5+gxZ8SNBrhj7CPDd+kdn+esJumXgF13cPaLBtLL8hhWzcaOthVgrCEOq0+gzsEkeykOEfDt
pNlq2AT/4p3Siylry0WGmb22cSGxFWkFMeFa8w+FQ8U9UIIUtSa172ass5ACVkHqUeXfEb12z/9u
j63CoMWP8sF5SfGmad8i+vMisaA1W2L917zsKXCgogUPAeKRjF0RzdYoLj0JVfL/D1H2jnP6bxMs
VP4i9x38IupEBsHoo4g2+gHQbOSwA036kY2+5/t5IoyG9UAioaujLikEWxdvvpQIY8Lfra9WIOR3
14X+4cNNvJ4k3BBONDkFbtaB/LmoZWiabLcr60Ki310iP0E3FTvC7x/SU1C0S15n2zhecPiZamSf
EY98FVkxs6U1Lgaqnl9fmi6infd+nCezP3mDSxRWFh3XXvOR8IAeahSy4ItB5z6mIZNtJyMVCaOW
lRiWjKV+f/gNl/H+wT2eCw4fg1AZTaczHpll3Lo3tx3/BfapBDZ+tMI24N+dxfTF7DWkm9dqBhPt
M2GRuSq9t6+4URdg61G14/mBMNEFT/ZHmkGP2ufzoWDUuXdlB2mlS3gGLKmn4QZ91anCo5y13VKy
tPXXv0QA30gcu+SQaLUZ9heobUQ4P3+g3V1YEia5C6re4kPCLZCu1OqqtXvtmUaVCzg9A9Fe8GqQ
EwmXJOoDfqgeU/OkWWZIrEkbFUZXBMo9ENuBXA0EU+MbmYeMQscjSxy3D44IQVmbogQu30C5Twd/
vPs5JikrQkwo0ULheIiDd0KdBDGs+yqFkVFoDKQpZmLv3q8Xo2j7ubieFEyvNqBgIUSbBBHLxRXw
CnSUpQ+MVXjp1O3EtFOhLHuH8jpVbAUY+2RQVhqiPBBMdxz/EzghQBeov3JnKr6zN+1oRkKC70TS
kBVRIGBPHC0aJygt+Gy5fjqBaKzmYVfz+K7H1Dai/MTQ08xsXcavRsY8ucfQ0aTaQhvi979gioHU
jUr8nSG//ogvMZjkI1tR/dHAQKiliGsXvz6A7MTo98MkqrV9ssoXK/WQc6LSE17+IgwQqTbPfjY8
Ww/+3MNbEOzMymsDJURx7wxUI91y2587QNaDleKS9BOevXLQsQH5vtsJIazoFsXvWW9s6iCW28Ph
umhMdPnwFm6FFaUBgWoFjRUZItV9Cszg4ZqVAWNfWm8FRLK7VoEzsbFtoaOT69lO4IxwmCKEUBdV
yG4ASVe0U04cqpUR7zmtJ4S78+U25zMObgoQi0o5Omz/LOWfG0ZslTncYdQbE+7slfhMq5a2+3Et
rxemHTExzfoRDu2ndlnPgJ65+SlXoTA3xJMMimXO2AbdLlf/FAShMhiNo7akRN6Fy6wSFhWz3sFx
gQbOsfVdyYPM+iYm7L7cKw+wOHfHTKuKjZ/GeOBjrZ/R2SCrd/rY501JWl8KELHBB76/IjetY0Bb
tIU+LQyMcJjQpPKATBW0I2Nty9ADXGbSo1hV+je9dyf9F7QPvXySwRzPI/gEwAOxbR/Ckm37WtLX
8plTfIlyoWpjIpMOKMyEC+NxLSTupdYILN6LEbkxa/5ddOlCWsJc5wdaK5lRsfVGD9WbU8u5pavV
iEhkn19EQL+RNx+G8s13s+OapcxaGJrDntLAwf03P/maudBpiT7+QNRJHIOGFOOKo72S49AAR835
mM5/WeWgddn0juYi3M2q+JjvkwiB1vWyohGb04i+yN0sPy4Cu1Jv2m1+m1yUGe/mFAoA7jWUgiaA
N/hpz4n1FkH1wU/SKwleorFGvbEdl62RPM+GAU8Sey6AK8fvXXAHAmQex50s/ZaytN4ggmSJqc8E
2uhjYzHvw85dXyi/cW2oMtF91tq/5jzAxXguBtjUqjaAzZTPWNNZvAqKDwyYOcADQMB5g7FQDIjM
Nw2iSCFECSdbcO1qjHmdMSKm6e/hvYW54333i+CoI1tdyT8bxLu5AujX0zXIRVxsrV1104Q1ez2O
fjxkkPQlJMEIC5jsglILvKqSdgT406Ddag1HzPkhy+9hz2I6rrvvkVSZkIzD3gWv9q2/CylGEaSS
utvuE6Yxjej83rXRWoCVuhPBK8adHE6QdzRCr8IgLdJR82XbYrTacJugTqs4Fuv79YvE6xPBGVqO
y+vaytJtSfMO2nsL1j16h8jRNZXx3cwPVHDZlM641i4hG0rBkOxhZGGihU/Ckk1/whRf29Xd4cJK
sFVVolahoosmxRAXmriyXdx4o4ARK+17HMUDKeK2cZHlvaZnVcDOn8U/ihMueiPT1ThKd04TolqF
7F8440fdiA/YmS1CoMRK4d+hJOs6jsK3VF44E8TtWp1dEYndbukBjHm44lcfMnf6f2Suifv+rsXV
peRmCt1p5llOUb4Vnuiml36JpaHPqWUJLNMn+zhLkURBJYbwHYLitoJXgzJFKWsxavSefGkbsMZB
WqAA86QjxnI0tH5PbVQIdW9Tm4mP/Ut6jage+bUftW0rMvfyMquztOmsEIa56LtSPE3AoTmoxMQU
kyTJdwTxAd7DNvFOdLiTfcGFAq2pXA23l+J3Ug99SDAFGSwxTjWiqyXxZzoYmnP6HUCXyjzvHJc8
PbOYDkzofQA8UrFJZrEsF1zzXVERfaypOE76u/fEpiBtTDjh2OBNAb8/kByq6GB3Jb3v1WOxjKTy
oSIQt3/D4Oiv13Dn4wPziF0zZPHzzBXZn+CuPWuT9b5xk9NOjW/zwfNSwGCXm8+NFHIBYXj4Eqyx
qZ+v2bKyohvdAXoWWVRI+NLlNnmrW/Q1ieLSe6G8Uq6JdDfcrhlPElTvggFLSoceZrUvCbsHa3xT
CONCLDQnvCB0wuPnYROJcGH5QiECzyCsKJZ/yacllNkhg8rOhVDCQBbrOstwr20RSHUReUPdcf1w
lZVv47KyRoJg//AY7U67uSHQHV+gE+RLYtZuiOGzOodJfH+5D8N2V/QW8zjdCHYm5lxkdqwpRsyL
K1Da9tgI2DyxgtP82PMeI2FyHGrpsSNfQJb9A8SSfFdWuEdbnspjSWQeFw1F2T/wLmVJhTnVs6J+
5Ka7gzDJ367fO3SDTJTwX/zmAO56a8BRHTow7f03HzXZD7cHC2TGu1ttYYd6yugjmrDeS/6RHsc7
hE5c1f5HYjUlprHIxFp/ivim8bmpJfqgVeA8XwkXjiaVP4MZR2JqPPvvG1SCFjF/UFojDwxG+k7+
yhCFEaGnyLGpETEk30pIYMc2M2WOLwtngNtVFL0KmBhVhxNooh17RfKLx8X+lxIKvFm2hlHYFW6g
ljGCLlaD51dqNrr9X6FiKhpueFF6cxJFsSNmANZVvXPQvYznvWp6IP64xdZxNxHh0xIcBkILv9ZZ
nQbNf0c7yv871XAa3/i1pLklSBnq7RrTCG783B7NIyBD5289nvLM0apXvdjojKRNuhi+DiQoB1Tx
jZk4QWeFmVt502abM9RwdJLvxvZiJKIrQVzOGPtZbqcWTRYLfcG7D1xqepMTuo8DC/RQD76wO+HW
dM3nByyGds+Hdt2a4BRFZdOOskEaR6Z4h6Aj7QkZkdYd7BluxLhQdbL/zZ4J62NQzUzn9zOunc57
3gDgqJu9dKfSNTjjzYDTNmontT9DN1xxf9wX3whigffRqTPu7rISFgEKtmwLFQkS0u6+/Z0Gb8Uo
yw0xzXEMJLRmEzyDXjLdNOAp9PVRwz4Z0gsx9kQjpvjGIgGfDoKBpVbYEi7Jqr0hGzI7m3UXSnfX
T2QNg0II2fzmAyWqMxSKnVnOorD/D6COP2XVqSAUr3nLzFgrnqdpGjjg9SaKuWV3cymK89xuopAt
jpD0sj1xHsFKbcHOXh+S2u1r87Kc0ieXCr4OiPWymw+iE1Etsxj8DXs7nejZGUOz8zcPfcVdwJQZ
o8NtSE/aaX5dxMKr2ZHMm0okK/GFYMfVx9q2r+evImDlt3I/lgwO8zg8BclBhPnwte1qk00mNfO2
OtJWe4xW1tk1K9NRaFTnpxWE92wLtWjX/cY3tcj7vWI6HnlR9KEoFp9AWThVJzmPMimzhd7CddAj
GajxDyx81ztGVil7caLk3+edurRYlmObHyHJXFVNJnzU4QqaX+n6MvH+TXaYuu/gyicJfWyoP+I/
g7MRpDRoVsw4Qwjuq0T9XP4EXJPNt0SJEozNLLQ9RUX/cZcqUhkfay3Xj8f9KwgNcSs/JQEQqgNL
Wt+FcT767RLHXbWpzyStn/uNbSGoYy5J2U8/qWStf5myZTqvulVOK+gyEWh+fYhuuF0qCfZhYl7d
3YjZ+jXmTQWmgfEVV48zYAdEelPTRzz+TNf/pCmMmMg1lwfQIlOV7OiDe5KyyrfIQikiNtPyv4O3
s8T7jd9JGQ0gk/X8ohMWODYycNXjtDn4fPiqADAaP9m11oGE7G0U0/+EG3LbEG8txt/0NqI2+pdB
mGlpFbB9UJO7EVjVzDjQVDVchSDX8rC5qNpp5oIsIjafo8xAAAmvLrBMInzeJmO9PANlyfi5b1d+
v1MB6UkbrngQezZBbKrZzXg6jejhf+llDjNzUSEkRPXqfU9f3lrQ0z36EjByQ+S/hEkd98uUCsIT
qiBDvg2+/YzmWfri+JSm+kU/hCtJZKi58jpYhs8+/NVY7BzGF2F2pz9mK8wiRILyYjoEz6E3sg5Q
Edq8NUjdVXABkcxlfcdfTfFg2VhJWyNd/HVEorddHHD3VFUpK/E5aYV2CSmYd/4C7XKqOMDGXW81
c5MW8H9BKLa+d1FMMTxnfMRD5B0tOiAikalmF0BH3Ln6GScz1xT+8oXSioJYQmkyYeAOKmFCgtiY
bg+xHyG53tJ3RZXrEYiktPFTszBQnWL2h5VrR8Aq0GY3gCKzCzOKCU7itpKfngbQfqEe3kG8CeOF
jcUaRKBf/sXYSgNsRog9Nc0UUCaDEkOAhVOQVGHFnevUgxpSVxx80Sb5lF3Gj5CN9K4BFL+I5BVN
NORZzljjYwRQOgVC7oeVRGhR1HR3ydBPhbjPBHUEdQUHrKienkN7DxAqds8wwrhTXCxCnhovNrOM
QfjhPpf9PsMXx3Og+AiPKDTTbQotNaJFS6y4pPE5NVsi79f+/RXBSVfKry87/lUgudKezOH999gm
BQ8S1HYq8QvYs1lTMa+CnHVz2mPy6I0LBATAI+RYHf6ATFW3DBZLaNs0/DcpitKo6RZVgwKY6u6X
WgHiB7Nq5Z0QiL90Xx/J0r5JLerVosgo+ShDvwUBUT362BsJhvygMhBB+hFzfjwrPM/BXJVAlA85
uvL2iDKzdikNzuoGSlimBnOkUhtjfu+h3jo3rZZj3w1setAQoZWlVDJRbVm7Mxcnm2by5FtXa+Hc
qqYPURphs4xvy3CVfd+ma1A7ZBWl2ea6a6GjPZPzVRRYYME0T2qEx0iwRbQX4JkQuArrc6RELfrU
etTmCwHHjpDwlT1mmNa+/4NxoRbFMNldM2Rv5BcH5lsBr/ZC4saKTG5ow/t9yrNmPPFwwRQTL6zS
We4uECpiT+SKoO3qmIPnlTbmieQOlVGTNX10U6s8SxYhLU32FosF3DnW4BGyejFzNNb7loeZ1b+K
SWTT8kBo0qkTS785u2kVE69eF5nlygdxD0k5fuJNNxy9F2/IYSDO5nkaYQI/kDeThYiIapbAyWQo
1nIumiSoKifj9ppMPJsoQjDIVSjhwlZRy9JcBCM/Ob7rvQsEpgUth8yzQye8KK2UK1m0alraYSWk
k9+s6Kd4sTuY6ni7o0zpR4WcP+PitN0CLDT+sb6diKHmoHvhP9ccuy+jQD+hcCi2Vr+qSL/U+rSX
GDDHkAOm+gn4lVC0yW7cq8tAGQ2zK/krFjqG1rDu2YRVilLIFjGmZcMspyOlGW1A/42GWcootsGx
FHWU8nHu5UyUNwaHPhgVI0kLWZkJ9jeLwMiKC+Y0pA87MnsxOpmX+i01no7/Eb98bKuwwgOsXOUo
9lkKQ+IycbIcF4zghkK5R2mbkwdMClePcHi0SNQdkgRXsDbVUWPbVedo1KyULZ7mAlTlHAJvoEoD
oohIjHfulQ4WSngu0QTBHa8TZS2nIXyvVy7hSLcmcxKSkfl20dafOtRvZAbjcKczQj7REZbOTlC7
IO4pToJrfhWxVxpDHAZe8xd/uylzBfxCAYkuvFFt+r7228a8+hzcz054T2QMsQFPNvORAdvkOVM9
Ts39+0GOzQvEsmawTnn8SwIo4B3TzZZRwkaGdbhX0K9cXhjvzmg/WBbn6RcC4Irx53GdLB8iJt1Z
XWvMBvgaxnrjCGNjKaVj35wIJ99DbvzPPcQz/XhMlgR3XBqgezKDSTbBRAX5v64pH7U1KUvhlohj
c/DYkiaZL5Oc1dQbB553j29Wtuwv35hGXiNu/HDQEW8B5ygJSoTpQk867PAZudsPBKZZJQsWmk3c
fyf+VK68z8LP302cnr3a7ldKox5jJktN8mw2iEMw1zJ0sE8oZ7vdsNc4yC8rmeFV6jbY9UiqeRmF
urBSoNeOe+WH2jv/vAayRRD1KUiWTlmjq4pBWldxkNJL4CFbH2nTQGFLVwRr/W5ydMUiSF5Y8fOK
RV/aJm8SEt6jkMD7tfwyNLngpFGlpDh7OOoDy8Tyq8ODx1AiskRQtusMFAncOVq8oauVF/CdZHtU
LlsW1awWmT5kfXqSWEqk3vT8qIHia9v5FNbE3EuIrshSBnhY1Q5QwkP1v1ZFAF5ErAozLMePxX4+
WvevvPSOyNicLJWvEQfO017HmVOUqtqiD53GFCQ+9UAycZoUfpgD4Fi4dG1yYZq/sSV/hodcJQEm
QBdRC2oqnr/Zpb93odqMHKSysqDalLOx3HxECOnMHr+CuLJF2gIvAFkG0ougj0JaSqklDbLRmqqj
SOQOA9VNY7wScyLTrR8ozvflvAa/jJKgDDHtK4PIuJrYQmJqUlKuxadDcgBm22OMQYhkKOB7fluV
EgU8QxsiGI0QFP+tf43V/h2I+2kk66RNYFY4lfavhAkBkUn1JGngBndRlsWtIpWlwL2z/NIU/DvQ
89ct1USbyN/ZIkTo9EhUD53vsZYw8lODFy1jKVjhPhu/mx+Ifkiv7kN74PqNjL8/VIqTlYK6wKEB
jS7JlGgdqc7wkQ2gbx7bBhPBlqIM/Fnx8g+kuuKdMxyjS+LdhetLKb6+sDKNe/PjpBjBTkpiDzrd
iZ2L6y+PtwSQuJo2PP6KE9fLrKLzAhkOgPG6lv2+0Zr7bK/WvAuB6Awe6vdweErGHQcEA09zsBID
YVOpuUzX32r7SDh7FzBHi7FMumZFUT99pxS2xbq7zp0ExxqJSl1BY57dVvLETONDzY7xnaKA7IdP
GrGGL0/1HVKf+21rQ93PA+JrGufUnUBxBy84hcayxO5saa9jXrmPo4yhug1JR6PB8lMNNdZDwGTi
mf0Q/WhNPTr+R5uikmE+OrvaaAg8vp/pK8BT1mTzO2uG4LqcQQWFae/Wn2YzMKXtorbaZJpO0Exy
TseYY+W2VJsuTRMpuqBubyqsxyPtyUY8kLZSVmgrlVtoYPdC6YMjn15MaXEMZDtFtk34ycDK3Tka
7gYFnhiJLRxB+OHTo0bhvZPgSKzIp3e4Oa9EYWgbSmHcDWQpJuEfF+xfi4CkoZ1qzjQtxG7HtP1X
rlZM5uuSvkG6/K8Jar62nWLx132Kv5squQLQpvxA8BiFUf4WoiEK/WZHJjjo0+5Pk9U4bl9gKUjF
zjIEwnNWNlCBRaGOILScKtpVWQ8uVhuvjonXrIfcSrxu1J93BQBuvtf3HLRBbEKDoElZyc91rl0d
+FnzdqYIb/ZGKLRrzAfb2fdDvu9uigRAP70NpDsCcgTIQ1tJrdNCf5VAnFvfHnJodKDBOD0o/0EX
80kze+u9Y++G1w+iUYf8ytB/fyolQfj8LPM+rZzKT8Zso/V6ii9PitU5rlO0Ef9A1iiqaEZdF1JU
hhMfagNsWrT+J5al/Y0PQjOcsOnpyyQIZ+0q567kplD6q3AgIh/p87ygDift9p93tPCjd/hI7hV1
Xvd+RdeAYJN06zmOdowSNwstYU+vQNPF6TpEGCBB5TkmFqKj1irXkDVvi57HmT6bH1z0x38cl8W4
dZl+KSbMKpNPBbS/L0cE5L/a6GXVWr00mhUyUGI8+vU6HmnGFi1mtvd/e56eZaFH6zSaQDmRWYD6
VL4AtJjapcsob9t+tAj+WmGaXwiwyi+sDS/xdT+3m7dZxGCk9fqfZHosecZkkAD9SHHbTXKonE+P
WXLP2291lBB7Ph6KMRQPEWPK7prOuAfwIJoZMhIvEbHuTUL44OvpL+6VA6oLPJqiBK+PxcDP4I1e
feYfAxN4Cq/WpzP7vu3Dqx6lLeillkIFHBKtlpIkdn/aRScyz5X01wjgnBmx3IzN1PE65uKfAiZn
zv+ZFXrEocAzNMTC4xNI04ipujBix0H/RLUvtAsM1Q7Keaag7TeenxFsrv/8nI7R/i1gEiLHqi8z
ixu7GwaHqRv0QcVpN+1OUyzlp9qFU/WSwFj0EJOfezbG45G7REN18MmF43Y7JABC1fVMe16jiTBY
ZfWFUgze44azzV0nC42prfjKP9lgSr0VJZzOIN4s1DifdH8sqXewLnzzW9s7VB29EGWCzjvpCWdX
zeSisc78MynKWZ4T49OuF1NTk8KRjDCRmjXGlHKh18znxwNxqtKjfJv9If8CO26Ls3/j+/QbK6co
VxRUv+FjmqyVpCr70vVjQeLa+jg+xe85m08oaE4pOZ1O0ui4t8ErrX2FjLAG1+v1x33ywvdWeAlP
JMIcs8sc7OQPPynm5nLo3rn9sdtfUSxYutWL6bZsynz+NDHOsr3E8Koar8t12fQXNLjt5RdAiBUO
cNPKGHvUYthJ4grTEj6sbCnLafv7C65igRVPtnvlhwAqut13vBJ6XYVyxHg16pobw56GohC/CKDw
1oZTZeEVn+7PnK38UFHBz0D6K/y9KPJUQBydKfC2l9q7pBmY5LbBLoyZXuelHV5I45y/ZUW6xz6j
5LHl2+1NqTl1DeDL8OCmad3GyF8ODhqhZr0ViFf65ictKL9d4L7s10UAAPSwk8eaDL0Yu1VVwZom
aVc/ds8aOreJn0dG7+mo32PBMZx2miTkL9edyQBIl4Zc/nJfbZpO/VhQ62Qid63cTODFwS4FmYuR
Pklcz4OtaxMjrKazwoptpu1XUN8SN7pI/vHiXygnfp4laTjB7k8nRbP71x5VElEunfFNv3bJDxWe
cdMEvUqq4GR6tps/xIyeUQuae011/pC5CS7OniGhWDaWHruFOzwEHNW0A+pJ/yp5CNLcgxWps7m+
seMD1OooFvthOdpuOGEgGeP8UlbOoAJKzxgaJuY7BMrxrN4cIC2d5eASr103isd6QHZdvcB7bdE6
ul/elmccKEf0v6i7PfXtC6DlrEQY7Z9ZjpoKUr98h2iUza8pT8+oK/jx7bEnNwciQc4qzCsc3m0b
C32ABkmGvW91c7Vw153KdvdN8kSUN2NZCDjmq3ALN+XUK8ap9rkEZZ1nikdt/hxowsEj9vOBxTg+
5vWRrQ1JfzVl3gP9U6SRE15Vb2wCz9QjTHgzI24oTQYOQdVedkOnY6QhB0v+Ir3KtLdo1sb7aTfF
NN5YLkR5kmU/gPGRAaX12hjJF7meFQ1ACeOLi0npCV4fy0ciKqqs0PQK6iRNdfrbRB0haXnY8BcB
PCSYnAGLvIE+rjtdNWKgXmAC3vnJg5HkYQv3Lj3KWfZGU3N/KiX5EF+AtVCtYzcX/y8cFjJEGRuP
OnwwtBmiAhmZbUdkIjyU7WmMMQgw5YMHsEFUyjpjbh6+YyyK4R3yz1O9dnTcpVURX24BdXKeZPaA
4/su/+XSdZhEA+ZHnQce2Y0Tj7WbGaLrHaKIpcBfYqhNx8o01/C3HOSva+6LfWiOBWHv/SXoIT71
DFoEEcSz+hiZ5QwsAOs4eqZzKj6HIPgx7hoA2latqovxVifx87H09sZmd7s8UQUT/DGLciK3vVtP
lLuNqNbnx8pAIHJuZz3TPWg7MrGnYNVsBkgo2htIQeHSwGP+2DirfvE1VZ5CUzlydfP8LH2lXrWt
teSagxSTt/yWVvr2D/MHCS/Qt0GXXja7GEAdbEKQVENoP0sYw4I1dQ+A19S3bmgqau93YHsKaCbl
/6u1J7B3MdLZN8TJxoP81dYzb2JbfDzS7mBXzj2hLbJQBnRU+zmn1CLKjfAd8HfTfKbG3UJ+/e/K
xq5c/F9hPvbyY/39DAGGGImVv1FZEJPXon7E/SXDUSbsrwlOZf8nxIduaQNCSV0BQ67ObhjrsnEQ
bGyKb4uTq+pIaWcaeg67QEZDumcmki+/h/amFOIDS9hA8w8ZkzWA/MnaCMxPG6QvpE356bP8qrfL
HR66658z9PaI/bIdWckx5QptHflRwB3Tf7Qsb+u0ghckewwXu/4vtOTUQq4AMsi2pKDdUfBtAND4
5KWdbfaU1g4yU4Gr8y0bYkLKMZiuriqkqnCEMwMzeWlh5XwxW3Z/z5UW08iY57n6gWmoc06hZk4H
mFvv1G9pnCHVRdNxe+N30OaEsYkHD3WgFcDY8xuNn0qSXiuKwn87ouTodLnaFgc9OjHtNvnilt2E
NGId8jDQB/ZS5c0VUrMnP7AwsjZ3tpHcToZ4gNo1Lx/OHI9iJrHVJBX6ul7xjOl7TKYIPps1q+bI
FXLSXYIbrjtG1ttG2/xWHTF3+el6/1elCTFQxH+m7OUI2R+hbeTtOKxfBcybNqqeSioXgb2wIrqs
tGiexAo9g2dClmK3F4SDbkTfn7w+EqkHrxLHn3AcfuQuXPCOeyMhRMJWjgNzB3OvphZgY59FDwAZ
iTQc3yPSZHfYWXkTGkNOIebwNo/5TrnLlwxhgaORG1aDLp8Tzee5ECQB1KVfLamVah+AaNaoDYxn
WhxeBzQb4vR9tjD1z+iJHghfT6WMeYaxOygHTx4+oiER182YbJ0MQaGMcR21Zbqw8nAUlm5FG9sG
ahmoOkfKFoqPpVsp07u+RVYWj1wvzbQmJW1sXvyc5tixHM77gYUFie4SahS/QinRdTINdIZhRsBh
uJdUGOYcB/ZEc9+ZuoD8wKE5hGVNNa7aYNZIExYGOGrl0V+qzz/XFtxfEuo1MpTeGs5vlt1JrUMq
gadAj3SgvIRTNJJFeOWg29wHUshd4YOTZsrv9T5diC861YLZT5+NQ3IsDk+rOZKLwKKN4XF59n57
hnoJSpH/UVtG/aJTkPOZv1p/lyod7MEd1Ymx0uupySZ1ohFGQ34Y2NEJGVA/c3FvnilC+6Ew/OQN
n9UymKlx7uL+wkW+e5nb2wvWpV36In/u9QvDH2QK2Z1wMUc76XZuD4OnSSV87lCEDHnIG0v2mmEd
Q21WSdqloySVSMIe84YIOJECVTGQ7qlbpwVQ0MKAnJESDT3QUfM170CKQSumrQ4c4QtdSlQ728CW
NgNBNCESwn/C2MI62oZK2ZRzAgD58XS9dxpeZkxeUv2YszvNiQ1DPdluZYlgP10LYsgCtFevIwsZ
tWxEq8uxEakE09tGqyxaLNAPjpDAqsL2PW+9nP1y3bBj3PTgJ0bVk6wDDDvOKBjkdYmNFBp2qm2Y
6DIGj+vvIlsTPClNH0w1HmDb5kMyQOuVYLR20yr6d3Ekf0uc1/AlmlGXskPr9E5Zz1NILPKZ3hjV
P1s0RDjvIdqDmu290msudHKb7dZk2RKedahosJpXhJw+bYDkuWJy5ecKHzWtugN8l0aKLApVdPhK
m3dS1Fe8BAMfA1Rq/Q6iVZ3HPfHij8NitULna24f80HQITU/V6x0NKswcu0wFDAxBYVw3uVex5vr
REtkmqmmCbpM3P1h9VuMHn2E0tW9HNqeh2/Vmra+jQdNjh2nd+c4x98q4Rm5ptuO36xKCflcvm2e
eBlnGViwF48tjk7MkIAHwlDQN0XWJPdCnMpnL90NRrBIwf2LD2FaR4Iq2jvAzPeHYtZ4lHkWcZZx
7IWdm1NbfaqAcn0q46JVNnUNaHAQb1Fua/O6lzKapxx7MCf3AqlFmDZ0o+vRvnOfhZ7OlpujlwNO
Tqfwx/n2ZTJb853H6LPnU7oDJ65TkSzfxA85akRLYoP+eTi+ONh73C+ybgLihbDM7JcVjEA1/bMW
1uwEst2Au7pi5xu3/PvhVfUrAG28018cDXFRDp4PwkQ86Z/nAALRTWXObuGNMSf0gL+TL+iseJ23
yWFBTDZuy+jm/C8Tbare6BaUPViRKwcmTy0JrfvAv/H2zWzlKUuNYKOl/hXM4Mu1wOqYvRoMr0tf
hlM7sDH5z3ThKwoq6a0bBHNBLvlN+Gj6S+ha8ygoDkEvCQFJb/95EoeD5TBW0+KG6KK5+qQHNW0m
bPPZVFpbsTfDRF25xF+Y27B66+gv6e5cH3T51rzeILaoZUclBAd9uuD3TXubRA9y9LaVT/8PimbR
Cf3Bxl3s+X86aYdteQvgRwLsA3pCCy4BPqiLlCTrhnHh1XhaYUjQT4vbzoNZnfru7q0oOacJSP6u
gf2Bw+8sQSh3V245cIHY85ZMuK8gwiiOCDGUxWxjPyy1GLHWMLQUJFGjt5Wm0VVgvDa19v/SBLST
nwg/jeMeghSbI+gGIXPqa0mP82f7DvXXbFfQwOz7LgNcgrsjIVWTNQFAf7WjZjUgaVaLMaXTnPvx
1U5J8IzDRxSU4XUwbuG0V3ZuF+SMdLE0e2myQo7mjXH7cPC1r3xOOi055qJdzMCqQUP/VxFrsYM4
JfUVevMeJUL56VcYmAeTsGVNSsaerd39zxLx3zy0YmyfRngjh8uOlcMOlKNnSCCjHH3S55uK/wCB
5EmFe1gVGx1nwrC5eU9Ow6xneo3liGvCXRUpZ/3FWzdHnzjvKs2asdTJbj0EwrAwAO/igEilEbq6
2oR2glEErqEgcp1aTJDb3MXc7EyqvNYx0AvK9yzfO9/y4SSXI4sPGEdtimoeisN1P6e8cpozAa/p
cay/22Up6h8z9eEYnguy/RXZVc5jyQrSU6dG+f/QS/1Y6SacjBmGI6lsyjJDOQ5eeer5OaApinGu
FavLEqWmm/y/fPwLYjw43UUiv9ItLGTodAynjfUyNpAiFzSKtlMaQUk2f2ibXwHeby6gqzCXOatH
43WX2X9PqI832mUR9k4MkVxQBAAlRhOjWxiU0knnpH9pJnoWU7ih4zDPs8ZYHo2Ot4dzEpYngl4s
B6CjHjf2XbAtf1Nm92nLy4Za4xJb/4+ps/2pz8/gf2yFnQoncCJExWwT4G/NlUVoBrOAo9hieHP9
umLZlYr4dnHq1gP4zfNaXu6LiYR8KHE+bxy4zmdmtn635uqXckLZrHh4hVvKrWAinFk9gjLMKlzg
FW0lWMBoy030IxmtyY7ZidsJofoIJCfDL3tsQeiy7MIVq3DlDKfR9goPMj6PpukdxM5yrcCFMHid
6M+vVfw4ukkmPcVi3s0dBAaJrdMUTZmk8NAa4b7J/H8XylWXRUysyLDDV5eCla448DENnt5BAXxq
fCb/ys7BDS9SE44ieDatLdzcWPvEERQlukCE9gm0YU+Z1awbx0d28ForUTciLm3HkVWNmJM/GiCw
x0yj07qXBK89qqtP4wZ3DfPGmEKctfBpIJ0XLrpAP3XD4OXWNIAMsh9k9wx1g9KsWLGDTrgZAEaG
837dVVpXCOccdV+WmTMgaRI0W/RdQTab3Maajy2pgeqxMCowwPQpMFhP/inrdfnfYKVh8vh5sPtC
8DjZu1ovMJzi1yijLjM5gnJMZekCqR8oIK3AcbX1fhyBYTuNeK4DOc2oYXAhVbDzG0uSB3gNVKst
bjxCbw7aMKF6bnss4x48AJooZKchqoDpVt6XPcuzIohB6NeCakwymeN9jiwaywZNp52hv1z54akf
rfLJM9AV/ybp0efPSyVVKDTfsBZLerQfdPc5rb97dtgV6KoMFkzbZ+OjAsASwn4GTDu9TTlA9JmU
TgT0XfvQFMfqvbCnX3eoPMgK0MQa2Gc5KENo6v2GERXvkSjEE1DuxuM943/P8knKkFivka3AHLyu
ryfSuKXeGvRkwqZpHBfWNJM6NoDxpyyn0NGkZ9pYkuB9TdqT1L1zt0GOqLO9Y2hM2zNU4zlv62eZ
NymE+rsNWLhKRVMyyAngJVB8DknqpeI4KrWe1iKuYi/iB/p6qcrQzyveIpY0D9dQRqnx2Zv9vOWQ
aS3XY23Pxo2YT2/qnEgLIxDrfNHnXenYtvZOXJwPf24BBSHvy+t23NnS5avYxbGn8Q5PRA2Wl9m2
R9olEGCbP5xxKwH39VptvUrBGWt1XAydx4OsfFm1A4d5JwFm7yikWObC61eeASWXROUzE1LAvtTk
05Vv3lCOMheJtSv0L1ewapaSBfKVnWTy/MmmgjH4n3IDm1zU5PH/NgrK1Npwjdc6aqwhZz2Y/tPI
7zR8n9zOl+VECYe5MszSJKLgp7TpxH5zmTl5dR34IyZFzUHeTkvE4+tqTOY21CLgvGCM47gPxFS/
mDzHFy6YDAcPcfTwXYi7Fu+Rk+WrwevC0ooc0s/hpGxy/a4sLnFZ1Vh1/vVY910GIXIuot/vp5nk
GOdOlIQeJTVlGHmo4V94KL4RUZ5mqpe1bNFlt910wk4mTN2lnkcpaBKMIcaggkTSPfG1p57EhM9y
BPBwWoHlu69TaXPumI5JqhFH2yA8GjgNOF77ov1BnvUQTGXmtQ668BA8dA6d34TmjzFf4qeUVtPR
pvd0Nzm9RMBcz706NlHILE3Xb2NjRrd6KOYgaXI07wewOcuX0T65nYMDwDL1bEqihehnV/veCxJm
O1b1C/Jqn9qC5Z/FB0jcsz8aJZiVHCeiNNMese5edmE8s8MBA4D9+OaqRwA7vW3o4/6Gd5f77lLj
3qq2v7VRp9V1NTnU1jwtekEx0qH4EBv9u5UpshJZ9Ie7e83jMYEyPTx4h3gQpyx83enrB2eERa/8
g9BiUTdNhfJGrMJgxEMm6WM7J3wg0zZxJGGonOXyzVxQS0D+Ijm8b5YqPmo8fRHAKvA+ry5Nn597
AzsmDSj2QntjmydJcE8LD5e3GM6oYjBZW6yMflbHiTYYke0f6vayfj9gff5idgMVFPRXPwgk4Mmv
BlokfmR6477Ui/GY+sttr8JFHy3iBy00eE7Hoa3eGfWp3e6as0Q30qx6V2xHs69I+TsPqIW7FFEV
xfwa2NJK1+tNetKFysrYQGBx70GKTPbbzeDkuAUiHwTzHH+cymjK9ikLGTZcp+ZFGj3BeV5uRtoI
gaw/39OhxYLo8UwVFZhbkKxDMaNPE8/KrEMyuMGllM7g1w2P3yvh786AJR7hSlPVoyk/mf0ilSpT
gYxFJOy8IxdrwUoT6UXV6LARst7LP8I6xAhL0P5/A1K5OCJ+ypkA93Whr3cH9PAHnkBiHnGZu/jY
mPs1jK9nbynz2t6klrLuv3waO0f8W51Bc9ptiiYAI2rL0oDoSxXYQdFd2wb+N1v7fPI+jbG7fkA8
OV2qj04DcdoxQO96Kwy3PtlOtgoPZalli7rC/0LAXsJJjZNbG0aTnpi72/VX7OuVq/KiD0+gxO+c
0rpWDyKcgLk1NbZ6W/6pJRZnNGEneDi6GLPBLOPiXAXt+dBdCYoXnFXWkVPkGqmPviTOODZLAJY4
MH1anI4y/3gtVSR/IP9yFkY1VIHUajKZma5sN4+IG47bE7SFUYECMl5hZB8klHbwTqeLOTOAXoQ2
r9jXRg5M/0EdX3jqu3Bznhfje7U9h6KwD6CXG1mM7p+Yh4ahqR663lot5bz1NfliUMlM1JFk3Hed
FiQyEFMc5dS158/0PifmFOZrFG9FMLRWPYd/GVRJZVRmHqs9a7/KgWW/a0f1qh/3emsa72aTo2rc
E8M9aERYk6kkfvWKDlV9eHfQpJEukdo+gExRmkeVLnKsi898CJ7Up2XPDfJalY+8JDUVAugQ8Mbz
cZK2jci6OiDAXT1LJjPGLdOYW67cGmxZxnBuTeddTcdMRsbCZ0l/O12WLKOQepZxfzG4TE2eSNwC
Q1NP1cNlD8SwtDcBCMGtn1j5xeCihGkqqicktzD0zxG4g3VQssw9OqwuR83+e8inRPvM82e5yoHq
EgqHm8dhwQepph515QHSCdcOc0hyK032WMLFF3D4bgyzzReMGlB7QTR7db4hkmL0EzZsf/xZzxhF
sK3TkCaQzDc4JE1MPb1IjVaxncI1ywIxXk+yQfLq4yzZtCkEQiljbPGE0cgcPbn28SJ+IzKj0JQG
f6isT5mrdSgXfIrQq0SP2mhhQhNTp6JLNNHDEtsWzP55RrtQhB1kCLgGqzQuL8Wg+KCG4o024E/N
sTAAicsLpUkcWfQM2UOe54YOZUDCv4Rk2sG7NSPpGKCI4BwUyJEgIE4I/Hbd7Hr7cpLCHN3DJuKs
2kWyUMHDKDFh6pWjChVZa9W4kDdM5u0vXnTW8pcKYvwRTlQdaZb372b9dIz6B5ezEd1NGHA801G3
1K6lvKNYDKXuK7Gg3tXmnqJU9JSbNQ7VARWws3rYJrPADT4tv8vLV/9chX0LjExTQq4V4uOYB/q/
VCSH6GAEnsht2Vk2nkZlqPCGT/RdR8vNSGVJ9reUCtLnNKviFs2ItK8AXhHDGkBB7e1Xsheg1GjV
BhIBWVtlYRPrBXoX0mOQmjMCQZsaRyWxvtaFAnIt8pHHyABSpT01DoKgiBI1goFP3ygxA1IfoaSF
wv7WgD/+U9/28w7GEHtzaAYWKZnhFfdLvq/zMERfCdnic20pR4/giZH7pIYEmipHWRNFF5sYSseJ
MaZpHIo0zkYV2tixGdJl1uFmqY7cOa6VB4QYOuOYO7x5JL98+JpYZJaWwZrSWmNMtOodY0k+UOzq
UBhSWyKwLSKw0sXKjmRjrIGxRudToPMh5tDvHWmjZ7Z1xAThFeBVs8x77c6jKlyzRsduJPhbCgUy
y+8SdosO+adBtkdO64nZXQeITZCDvmJxtJemqLTM74r9JhreQGRJkDfSXVfrW4ZsVl5Fk/P0W2V7
Ic1wQWsiL4cdHmNrXv3tJ001AVa021t4o6I6BVOWtc2TqnY8JS4zQpdMus9B12HPNg/DdTZlHCyr
pGahDLdiaRmNyJGC/fwKV7aQdkUnG/ucdDIa/mMrd7y8CaP4Hw3yDblXxkPJWGNUokZIcNxqaosu
+lqtGg835SGNlo5unq0uxd+1cZrmTKX+Fcd6TXsO+YwRsxYjNyo7CpWQG0ZG0A2hOSMZIDMR3/FK
8Ezj2PpcP1uOnGxH63yJ0CvJI6iYzTU3czTLdvztaleH642tJtVLpRxcMo56FlE7E7A75yQZpQch
pHnr4x/TisWoVefIc5IPzi6+Gxe5wBGn37kKS4CcN/tpj17lwrAQw3kVOyFUaeld55qi6eetsx/1
sipFctmx0+bQMdjWNVUDaURwvdkSC4tuktzTysEo2DcYePrYAO9pW+dSoiWB88JmwnlVovXkYIbh
IaPn+BmzMhErm/2K8V9xMUZMrluPBGgwIdAkweaYtuYIVubM5TxHWWnOdyGachK7kkD7sE8LPgD7
t2bILrXV9bwHmOuo/eycMzRabLq1lvOkiDGDdvDSbDZc55VHAE9u4rem2ZbjdTXdeQ3K9ljYQd/c
u+wYShC6PuFnSk7v1J/x+vbALmXTvHdlOwiuz0HkUnIPmBlFQ5suw9e5O8mAMYVWHiJyftvfQ6k/
xcc85MaoAUEEqNbVcYHtHnkgcTS+5eMUeKffVlkGdK34QB+A1D5RqTaS938p2RJD+GhtYqlNWzPa
nMAND+8eNiGFJQV+krbsVWPKuLEHz7bybd7u630s0RHJYKUrhQvFFt2LxXgVZ1d2/AWtwiu5WMse
ePhmpmwJbNyiqFrbr7/lR7kqyBkbl0zrDgK+6OYoFRaU8c+XFzI+CiooK7HdVZAEjeO3ZJ/sbbqs
hhWaRIruYB6dk2TDkHNvpSRWhprhb9o8YVe3+SH12c6TJVMpSCCjcl8LAExFfLbWFBgFLUsnByMG
v6nSGqKWMW6ndgsQc935870Mv9Uz23umlePoGPC/9gPv+wbQ27LXqM3NaNlWHwmF8p2xUTUPVtNt
5T25VXGgHebz7l+ENf3tSuDIrJJs3owocTA72ekWvCYBD2O/Nd50SSGQsUFj9jrqxMESD8yAXBuA
ZhrSB32KRyUqPM5d1VQueWeX51/QAEDjDJspvqCO6LKXB5lCtElzD7rMZ+0EknWOO21Ag8mYJoWh
iM5oGxp7HrLqX58Nuvn3QCP2T1g7xAoHL1ay+fI+GGzzcUKxX44yG2F/ztHryGHsWMTJbqh4BUrd
ustmnJSOLRQlN2Er5XjoasLagPzhpnwBnlcQLxSCy+xaIh3zPyUPXuN98ZzuZzBQ61OEvJuWVl32
bQ8TPMO3xdaeF+zf5dROlB1G2qjGAeUEX0FfyvxZrOoKawht4UvXM/YezYIA20sajfmrOA67GtW1
3A2sP6advHCfEHZ+EFrkqOaDkcAXpttK7cQaZyZPN9KyjsHtKHKxhwG0nvkP+ISH31jS9DojPgSB
NXnzmG9UkGBpyni3L6b6zsseCDV5prCYZwUVp6fYPsK5BDKKzRVI05vCspfsfmxSHWRjyREQI377
G/bfluc5BRcDDB9rGrBpcCGjOCZchRjkxxDUytpO6a5tkEOq9+Rp9NQxEG7PoVAYHKJf76FQWUg8
XjPO63HvQyOkIvqblNcUyPUvuWXXCGpvsu349rE7SZD0r3ahCteOrF8DYpwZfkCY2jGfCrrA7JM1
QbPaKeFKK0fh7Sw4xm4iSv5wbyJKwE1H0zkzIsQ21/xrUv2GdHBvkyRLlUAh5wv4l0SCSdQdVwFC
uC7cfIIZTr+d8PwjBuB0eaA8x3JbufkWYO9nQzDyzdaGriymLYbhJHimgbNkOMBhw5qM+w5ty5sQ
qXMgxu6grkvKDcBuz+1Vcdvi2JgxkGwepIF+USgqFxArgLUHrwTUjyfOZvD28RHuBPST2SpV9Su1
3CfpfFe3ay2MrPp8BfqgRa8cZYfDkMnWUkGIM2Odgpooj//lkTrIStKtFZnM8bUGM4y3TB08mSW3
h7gkSxhKBzXodVTEEpbIgok7wN/UgqEcltJ5watUTZkaq5rjE7Nrgs41J6JdI4Abv/VCKmgawq0B
0llVPF8moYLt05xUR7ayBl/eS5d0520YZvkeJsWaZIajnLi9tzfnL0N0Akjg8IjKRXHZmBj3YJNv
UGUttmaBc7VN9658i+OrDCmjbR6Y9afdtwpTpX/yjsrvb9VwllGd04p7himncmE0Cs7nygVWWbKl
W2piBc+HdLkPNJtwcEcBy1vhmixjeqpmBZimoHn1fpX910nHNzBWwsusFKwH93vgHpguZ8NUw1KM
7m8neVN+RoXwRREOS7JeNkJRp5d8Ci3W/xRIaWbVjcd7SKoMLcAEgjwlMkEYazkg2zC3Lj2v0/rp
L2ZIeZQOXBEaYiuk2YTWeyf8Eucy6dEoyoozZKM197BT5+dVgjLoqEJz/FtyR88F+qFAeMV68nvo
KFvaiWnH/VJNUie9fqMZXJ6jdDpND+RXi/tYVXZIdwJhbpUbRtlCydKWZCi7GH9Oo7edijTkVBd/
nstf1w0qEcEtnG0Lv6rhcEIPfEWeNPYINKeDjlvtRhPQbq6RMqaLTG9kPj0O+8cDmZiFlqVG3FAD
Er+KR3wtNGXg+qWKHn1TCWBjv39EgxAXwL8hsefJfbPnVr7txHe1ELQUY87mm8PlEgz7BzrqWXsU
YjNeuTjyDpf+dY0vckXlH5pbpDmqPyatX8Kqz5DMwhA5D84wa1w17hqO6MObF+6DXbJ1810SctUr
3olwu48MvfcE0PuEVhjTH101kUNmnomAqlJssbPEwG5nFlfF42qIrIvvMojsqAm6zZdm4fTxS4ms
ZWnFfuCSv7kc3UbZ0VN0zaU1lrr4Dw1fpF8+ioM2Ah6+QXLn/K/fTszNB+dA8YaQhDL1T8RFNZaT
Z6xSvOqwZtxV0RnZsrCKtkc72/e5tO+CnHb6mmnO5EBcHoqKilSB8EOuiU+ohuf4Q0k2JCehuGiU
Ir58eEV0OIwVkRY+DWAD6DTkmb0IibX6g2qyKK7+sinrDI5Zk/N4Ds4/KCBRiCVGRBDgpWkw3kLu
Cve29dXV26+6KFz0pcwZ5/JmoLLhKdfQOOGLTqALsFsbQYQxzcYRPdRTLcXItC4iPHbUnl+Fd8+6
wD5ksF8bacmtsTEBf+/kNy7qGNTg5QXspd6b97lD4YeEhjQn+Tfn8+ws3LM0smnmIA81ug9ZkEl8
WogKGlE+bXBIOPzjSiy36Aqix7GU8KWz0Izjs2YnmWX2f754FiQ3kv1I9uKhVM8USkT12eN313jP
5Xae96xk1GIZfPmFaGZwYJguPkhB7b7Rf0kY1WvgEnFtvhejiN1eyjEbOpQF6W5wwv0F/JqOicCe
Z2uhcI07sidJcG+Ad1w/y2RYYmjgQ+956nYcfzuzRDTEfQHZ/Rvefx14bfGNVIeRi2MeXMrXNz5y
yJ+/Gmwp2xWjsjuD+PhfxeuhjNH7Wu+Ov6G1aJOUQWyJthLn8S715ksXxJv1zXZKr1yG4n+0tjUa
yd/coSyWsg6QrtQChrYcHHA8whOr7VzU1grLkNTveXh9yjWlM+ueHlr2cYDfTbUw/JYgKiKhd6IW
kp/MAb0t7b1zaw0Q4RwaRnkH44J/kC6rWayFAZSvySaFzIkNddnzY3/0a3LdGsn8heu3eyj78BJ7
40xwUme338c/rYATbBiK3Axf1cwBm4S3suowLZcQteiyCCiciK8tSwQ/3OH1L+1zP+LZdqHZNVgj
giydP472GHuMH8rnMlSK1w6L47HCU93IUfWSwJ1n1cYFxBeYIGg8sdmrhGJmmEqbZ4/xosRfJ1NX
5trTIu6ll8MiGyXhP0zYQNRGwDjZActYvWZ0h8VSPajMgxwXMP5RYxi8LWdn+VQYYuHSoKppZpnY
4OINN4+Ov0kXdtWVYiMNJtYoV0lSt4FAmjM9fChYsMEuXJ7G8Oa0j0//bEf1uA1VhKGBcbZO7Kbf
wHmt19YxV4mUYitp/+jQRvH9DSnpiXp2jgB0PBuwt218YqqqrLvwJST6vnQ9mBqDxtcgvesDBzDL
VY/WCUxR5AQ+XLQdDvlmX9SPvwut47/2wffCYgzwB4FeNYXxnrdljJVeRRd/8orBOuLKW/NEd6d5
flNg0orXwYXsiF7NUibA1syOlpNTBAlONy6jUI3H9K/cC1B0m2syiu1QWDCaiO747yB0CUMfcLr7
rkHEA/bBiJ4yP7sE5xUHJbXNCdyTp2YTwXGzU2Izxaf+UxVfvu8rXnQnXjXl4Bt8kRIsqhbRLVQX
VyB11CAdqMsPyV6djMFbw61v7gxT3FEjlCbV1yl5llUGPKpedJ0rHHtDJ3r23Ui0cGUWgHymn5/S
79qu56Hgn15n8MypbSGWXxYek1L0zxIuzCG+qQlzBYelJz2HPR3OqNf5O/JOwJ4wVDQplrSGu1F2
9NXI1NbhXzFnWPB223fOAlCzZVJ9bBZotrnWyg3KrjC692dtDR65KGLOvqWN6vgR+KytoPgHtPRl
5rLZA2jPwrFIPTHaEZx34Ta5J1AIdud1/IShZL4/Ae1LWHtZoGBQ3ZX4OJWMkSrIELDeU01fo2qM
TrvqQpVjjCoWjBLcVxc8IOUqg0ejse5lzDFi8d3Z3wM6KmkA+EMjRHzAPDkM2AQyapy74Lnit1ht
nUXSe9WH5YbdruiPZds8i1l+GlK3R0RxAAHztKzGLXg+k121zJUOjr7LA7Ui78T8S5TGuh2cp4Ej
8Yzq948DYncElIGabFgwu536NHTIV+Afjql0yMBC/OUemgyrOwD6IwMnwk40L+uoeu8KL4nStC8S
aFD0KYSJAYJBC0WCRCki3rC6Mi45iiP0P8K8s75oSuxT+mUcn/yinJm2wrL3wpk8Hm+wumBeB9r9
Z4+Al5oJIjxIBuD122uIlU6pSBQbQCW2Bp6kGjQ/7FIu4SiMms4Zf2uZOgRKVhBDgNHTEhfPRhaZ
4dmWDVdpZggJHQK0Kygn1HyxQfTqwg82e2ykcvW6PhSvBR+bRuMvSoXLSb4exZw3zJgvBYw5hzv2
hNsqvkt7GntVcbobMKQWOUrUsqTUapnGyw8GR4jJtrGUppuMahaNqUEohR2Jcxg0WYm99HyUgdAb
VKdDd2rB1QGSsRkhU4zj0qiS17pubXQXOh3vsreWgbrA9g6RLmg50VVmvqeRPYLlj0wJudfqx9xX
9MX+Pzq0IsEwtsIe+Njr4X/QgiUbQJY07e0lSaVsKKQKWIGMUcrFq36hyF5qBasni/asgOG8VONm
lYRJg80Cbqof0l1e6L4Fa6tjCqF6TrRep+f8H8rtA6Dob2R9Td1sCweuvTE4i9lD40dt1nsJcJE+
6YY4+HqsQYng2UHKKfOBd9bZNZd4UxjP6Q1KQDSpn5yY1I9RqRLcWMAU2ZKPM36ekAyqWBQyHcaL
MRVOQiXIGFsBHutdO63Y4QaFAdBXyPlDf7h252qpdtzpnCgI1kTbZmNhZAu4teaPDcFynT3n9Rfv
RbIDeyN0lMIi3GaZK1b5chH24GqLElZNlZcA9R6Om9d9MGMAKoTwjjbxGJ1Mcqgtp7SGxJYt4bPp
LtNr4EM86+hYgKqWy3Swp4/RngSPEmWO4W+1Nc+VM81ze4HizSZj0OSPfDE7Ih6aCotit+QcM4SY
IlsGJezkLwsCgxeKCbnbvZtYweSPrTeHaxNr0Ts+1+W9nqi91CQMdWg5q00lgsqBAHCjCnqHENZo
zhAQaatVkvYNWiOOCvuwxHipRebC0SGvZSZY+tkZAyL7HrQBF44OdjUf8MMZyOAfjXoUGkFZzJX0
ZX6f/1aAzORdFzKk387Mn3XgsWmT3Sqgg+7u0M6+cLuSRTKOAu3+BoinArqb+xd4zAxrvx8Ckalt
PH54p2qs91Gs1FqOqQV8z2hRpoem5AELro5ev+qEwCnkW6usGBYZN6zna5ow9WlPsbUjeXHyUoML
O2mwU0ZI+CQDps6xephZrsYjMKNyeVSXG18Mnd+UZH6v+rbmTarbl6KiF5Krg9hkk8cJOTVIk2yc
Xbg+3+aBXnuByPkvTw10B3V7gMtm+Y6mAKL2fMM0DUjBL92SyAC51RO7Fmgzf/2bF9qcundkBj5M
yc2nnaYgDCctv14/0FbH4s3tuAWCDlbEgGQ/qF1wiLN2Xb9eQY8Sjn470Bt5bCF8MlkGE/IhgS10
jApohEOlsHggT5z6P07kiB9jk+KpcLHM7ns1N0PgF+6jyfLy5Iz6V8pChh0YR2mUXUudNvz1uTj8
FU1ldDftH+Drq/GgQxKE1NdONxEL3oX0fILIpx25eCUpTgnTtwS6mu/Sq5HTtW8OS9OXHK2m7+6U
OE3DVn7QFtOWXz2w4/xlo1Jg+PpOisqDi5xvKaVVlvlgrU83xgu8U4a65Mx+hwjnVT9YsdDtS6BB
8lMXg5rgoZIZ7bA3jZzCZxcOtrTepPkUbFMjMaFYK9EHKkquu2F+180dqJm0vBSUM7ZMrX9DE9K8
eMBPN631bKxzUHvXBw3va5CuWN+1EZTPWkL5QOfYIbsWumxPJneRHPYNYo8CmPXOZSqC256FXAM4
G6tQQgQdje+9FrWbJMlseeMFtGQwRLa+CW3SbmWxIRm6JxXMdRcJxHY8OMT73VUbwKXxRffeooVh
UP8xuEmYX/bAJ10GBe25PsrWd3Kk6If6Ofpb6BTMog/asfSHuiwDcnezJch81Uda+v8zLohaTUI/
jNeKpFQvpPejAaxBRwRKjE69oJmqsXGazlc/wu21f1tjkEAOUxnRiSup1JmnpCDPu8VOgsDilvsA
H42sBdXbHHoAm0qGzhavrj2UJ27jvG02AJSMtHXe5ZoHKaddT/QOPRmeBhznfGWJSSzIUVc+5oeg
jK+IG6ob76iSBgHkwg5BDM1AKQDYKZ2jTeCvf7IEMKY8gVCqN6nu+esxvFt+ksp3IzR5N3Qs/SbO
z5ugWpPHekkJZLuSsvCl2ANYbC//PvNYdKCLjE4Dmee/GNsRLwnFRdeJVZA/1jmEXimAEmP7zby1
3r0JVdgBkk1V019GzCT4dYTe3czeZOksepbhZBOyWy6I+2c1KISPiQsscEDiyboe5yhMZJ1VqE8c
P20DDOOmDrw9XdVP3APpbVi2BhklEVqP0l8rlSkMhRAE5GlZI+exa19+JQEwyms5FAIcgYQDM5q5
ZTZpjgfsRCAz8wweUByPfZjNMF2OjCQX8qu7+0/DSLmgE8/NSL84mNjr4Zn045Q4SXJu/AAsNrMN
tPHEV4GkPqG+AvE9Xnf8UfIeuP4fWysGdv6VX5NN5EwwDs2LrHby2J5adJscc8+nRHicDDRoTI82
FHcjldIHj3t2UFyuY0lN6poxijbl1o9Hl7PuNh/ZUDjionjoeuGF0J164/1YWKnTM7JwGx1/TbMg
KnBBQQ6pzKnTuq6e0xDQKN/IMu4gXJOk5ncy3rlhiwuUG9x+RSMhiPK/g/cCx39f1n/vJUSdvPsv
a9Oa9YFIG5lejUFK1/IZXbHR3hHit3CCkaYJafG7iIuVTHeNndkbKV07DoUyVvpqUiNcYwdhMD5E
saPbvA0wBN9gonAfFvBE1lbV/e6DZzn0usvFIz9OUuB99cyMqwwzwZIBQTu1KSCXRbLnBEZd+ovw
UueBsB+jxcJKvmyDdO8AkSaid5eO+/iEn3qfP1z+FAGTfh6QZGcg8mMgURj+Fb85oHKc2jrcJntv
xT0VOL1nvUOHT0gh2IYRXoNZU0UUxoWOVZJH4qXGXlFeZm0C9ZhqxRzFIG6nSqIeuL+Fkh58E41y
A18KSowcJH8PgRg+mjwTAS2DVA3LfYRVIAxflWZY6JAi7bVxPMySFkPxIrF7W4qbxh1hX0x7lqqo
qMJr6nP3kftthpxyT5Y0Ewdb2Zv1juIgYKgql8BBV2iSIbKAmkIf2Mkbge5ZBEau5OPNVsf4b7m9
X5B0w9aKNNg/aBTmjDm6OzCAZqkjMTBZesplPU8+5mXgjqZXZ67AV7hlqQapzUt8eCh8/bL28iQ6
ol8L2w7gY7XpllaMB9HoAHzPTpTgRdKK3xbdOoG+JufKMuUcl9+4xvCm8TvPz9yXGdSso1uLP6l1
XEs2xxVyWQ45JyqMd/46/I3YhWXODnO7xciWtWSs+6sw1Rw3eC/M8gLi8HfstsJUI+2aKF/vW4kl
aThChv0VT9wngoZlGUclCZ+lYYGhLI4A635QJ28/U7Xx0rBQ2r87A2QL2Zv1Px6LlWQsMTMFSnwo
ACiB1YV43MwpsduWljYtm4UhbIFxrc9b9mw2HZ+bay2DUCSpkc3x32gptVn65Co2xoxBmDZwXLEA
E5m4V5BvPuyYJtUuJD+iUIu1U73dnQ3+D9T11/YR24Qu7l8i4DYzbep6XJFtlx1No7+8jbVupbCr
t5MKO6ZnVdUcZZfZwVSQFvyzDn4otIzwpxCOwyKOrkLwryPArEEQoC5l8d+QP28gFCSCL2haoGBt
/MO+WEeUO8VB2EKR+U7RHS1fnTYUvtAJUm2OwkcQZLXDsJZO8+nd/oV58uttjxLLhP4tlE9cecyw
SYcjP5y7+B9zWPgmKnSzwODOtVJ9oUq5Smo00PkVAMFhLlCPvVtSWs2qcQCMYeviTHqPgRMpOMJm
xTa/T3vtL2E5TpyoRtk17zdWIZ265kSIYyIepILS3iXwbEFsqr3xxhpuNxYE/YTGrzRwN3Q0TD4x
r7SGOcoSLStXfQIbYOWvvMGxtjddKYBMTVvN1/yopu3sak/VsDBZr5F3UbQ/SHeDCMuc0khOW8SR
GD/0Y50qC6rAWkMODT4FWnesNhuJwq23wEMnhlxGCo8ISVRoRU5nIN6xyiBeCxqwWN5smNMgquEW
KB0ZH/dm4ydFd0dqrQtTS0HLuovXFa/0sWnZr2QgY0mkkfUy9NRxjYXMaIcTtCbnI37B2iYcU1Re
0l0GvvhuCvuyav6zo1vmtrV4J+N0EsIK3lFejvyZ6NXEIj7D7OIfANs1mdSui0CLbKsK6LHSxr6+
wKTwZsBnrsjcB6Yno5qrgykyg7m6NpJAXin+3OpV6xmxD7i0w5CMVRhBaLk5l1E8G1d5sH+PK+TF
Z1K6uxlqEbAlwKnJAIpthXt8kedyuYXs2oQGXbXkYzA6HiOXcT/l+XmbsI9V3me78h+Xbvok4GaT
VEz43y0o7b7MPGIHOCm8GZYATk8A6itqzT3h7c8YdRGk54zJwkfgw8NonDVe2TypPatQ5orXOaP8
+F1I4z7kR9VzyVYqtg/F+4ZwOsLg/7B+fC1TTzVROA31aQX1iB52DK1D8BfqkU2DUoB6Fkd4kM1D
qoa1X/Qh9pmc6bHY5EUpsCctv4citP8UTj/+TIQZ8IN+fE4S4w9YTLAXPRWv1v1MhkVxP+Pf3HfZ
iTFgdpjU/AIwKw78ar/r7fQv/BCtFc5qcltH3CWcnrLfDQiacI8vXOqvMy18MtaBs7zJ7+BTbnzd
4mDIT7hpzhD7xl5OaQ9H3Nj9tpGYSylArcDFBo40FNc3JBin8kDom8SNzVQUCmzWf9/EKmr7MBSm
EHCIi/USlJoeYEIFF3bP3JQ2b19CFmMaA5ZiHp4pbRTPfl8S9wEp65dZNLpFJIu1wgsOF48BmKXO
kxzN+z903lq6/GCy0P8pwVeASWw6A1Y7tfnya01/8HboI1aaMFDZe0w8EIuxWzTKZXKcNvzEE4nK
ahHbSV1OKS511ttbXWIQkIt4BJgd985zrY+GtHJb3+WfEYvpxem2E1tmmeRHPR9Diiq/VVY5s148
TiPLcoUQPyd8Lg+bAnLwzYPhKZTk63iYPX7YkS/h/iQ7vGoHVu1BZVQPOsBXUnYvEm8QR3Jvubh9
KJqspaHWvUDPY2x8Afr/PodrXgNzAHx8lx7i5BNpzX/oG82KglwHRHcVqn1rw98aY9zkdR5BPkgR
JtOyCSkwi416+KjMMxPc1UVAW9ht/Twf4XS2b6+coafixuEtI0I4wZ/y8cpdR4LqXAOVpCmv1QVT
nNRRPTuowTExOckYMK9+dyiU5PEvmqL5k5DWhgswgpBZPK4K4JZ2tYX56oS1VpnDdu80xyWlyQPS
rUqYf+TMFJx6MWmzp3B2wWQXeXLMqOoCVQq6Ax9Kx7HnhVrMCWixemuk/WBberPmGEog/cG/sGLv
cwoWnLn/sIHrB05OWiJLqod16RAJazgt44LYhVX6JeMlzlF3zmUtK86N+IRgNLrPhEieiLXRQtZv
0nxZrKg2pDnzRN5jlS4Qay3ZgLXJCjHC/Wi8007QWkKwV6JjD9/HYgTb0Wg8k6FjAVP/v/irt6RB
BGMBEIWU+SZOchNJtJR5wByxXuzoLPleSpFFg9Nep2CetNLg9Clmk046/5CKN71PFQ0DG3d6y5kg
AJgrDJKEwQ9yPxcXfTLtkA9Vmmgj0ewSCJFcAvEjuqSRkC4BtCfUo05x1JFLoq0qYwqcCQZAbORN
+rC8jlXRsOlkT3uFh0GBNCUJZcpb/nkl9KWRWJfBrh3agb5i457CjDxd9mjYcU9CuFAzoZEf/Mi0
oZTU8l25w3+ruhSBM7u8oVnzmq3fi6sLEOT7Lbb906wvrET5m+ZYdspTO5hXNnac24HIaUV4qvY1
JguM+KX/wzNhLxw87vH7/YRHm7fWdOUpkHI3X4Y9kx9KwGpIsFeSUWUB1tAG+X3yxpHXivM8rZMf
992HV5IoxuwMszG/k8xvqFjVcF5DkXn5Y1JG+/+zYAzv10ie2m2rcWO7UJ3NK3QFusCnUhsmObSB
Pw4RvbVDEuxvjsuXqQpLuHmlfY0J3gqammrWoWy7fhI0EtALEUEgWNqBYwduuwc9tjxL48JmimGp
4m8m5v/EIvrx9JsNeiae4twC3FkI4CXhqsS3Vz6PEiNdPAlFgO64VVsW6Zh9+pYULXFO7gJy0J2R
bhzVATlvpuRVJmcYvQbAdIKlnEKCLUzT2R+8HEuCgAKDpJQ7OHbFxTrwTVRUMLSqwf8Ipbpz90hs
ZoII1FjWWlDzF2yxfrdQWn3NRDgtkWvG3BMnSdoRuuHc+wTNMeuhcHLeziVBGZYorbYk0/ozYbpK
ZFLzeqHpSiE7MJonWsN8UvyTrf+6M5Eag34n4G8y4Ogj6kFTKjKCnYn1zQdOenknXHaggGNhY1hJ
EPjGyJ7XgbiMO+bQoKnyNiF9/8uwPTv2m70eOxhwG0rJtHL7g1Zr0+1/vG/azy1g6LqTudsG8qKs
66RnAoDVcZIY10CMkpA2q+luyd7YNWw3KoiUQcziUykY9ac+Val7Au6ll0i5cXhMDJKU5Hk+J8Jb
LvFtmAZW58NI6WdswdUpmPFC2D3/vdf062oBMT4o7DrhaXVrgeexBIIIfEgEzq1T0lzg3+U5bIfP
YFMow5MVahOguBp+glrlWm3khEFEtub/4mZL8zG5wZqum8wL1aeY566vQu3n3fOEa8O61WXzys/e
z74eRUm+6dJ5b3UrMlVlhJxWGn7heGbr87vA5mb3kzOFrWgsCAwMc/pUhPD9zSpWmjVoEXMeVhAc
qYh04qsNN2IGO4s+zizlfcqio0Tcqx5A0YYTWWZP+RW27L6CMsI6VW1uPVm3Fpyf/kpgSf0Ii7cj
I5u9cLQxaBUnyjHNWzEB2Hnpwp7Iikj2NcHH7uhPc84zpH9M7aeyPWiLu536lZTNQq0TaZXzMIX9
9fLPY/uDorldmwo+l86FNJW+dZoMw1e3ysc5H8XK7BgHEFoQk17+Q9V0yTqaWZuTW4tu/QkUAAkf
L2YGSCxGptcqCrqFd1HRojl9iaKFK5rZV5aO4czrmBFur+Ll2MWGLunm/86tZbdGQQ2L+LWnTnSp
4LyxEbtO370c7K/Ib3BlD2cE0Caj+x/J5aO49hB1KEu4gyo2CCUnKDghBrEN0LKOmdwwdSoaXcNO
HeGtCeulfKJgQ8rfNGcKLVOAYSnOiSPUBn99IfU7H3RF4QtP4uuZyw/fkTm1KX0R39oUqGyCrYEO
2touTUcsSh++CPVLp1s8CIkiBiLhwQvg25pUeR1ZfhGDzxPAn6YBG2yn4TrUMbNxpBh2taRs83H6
+VDUj78Yezp4sEDi6AbzH9D0UtDrz5G1gmP4lAYMzK9/qulAGBWgBATOq2bxx17RsKWJkbUNLt5B
AePDpv/2/0J2kbK7UbOOs4cvsltbR764vU4Ol+pIxjdpWcg5n+FvdngtuAvatOnrd49aGOuzkTKr
GuGja33lcimcGdpi88CwvOJngLYVhHBzx3/6G41Ue40VFMaRcJMc3Fg1jVKNEp3fiia1y0bthvzP
FqVyBicrsyLXDFKUzqJO7USrZ0RmauBrs8n4MVuMf+4FEu6raolN+QgJxd9teJXMs/K610PjBZdK
S7B6dE3IaGg1Gvt5RbUUo//lhJ/gNk/mtRvqoPTY+J5EBS+37UjseOh5x44ijbyYS/pkMGg+84Nv
kpqtIeeCb/Y6gdO7vHRCzN55CxBLIl9vO+1gT/zdH74g6/XIsxfw2yZ36FqB/w+7DTLWAhzbLNhw
w6vi4f/T/JBRORnz2XVtrrMTckYQji4u6wv6YjMk00xOu5+i9NG9tqu6fbcLsL8VhdYpYVwXfuQW
Rt01+YZj0P4yIY0ukJLvjNcgoW0KbwIJ8pFnCrdMM1dj7rVnoJXz6Y0dGKZI4MVXNZH3eeKjANaj
dsUFE8TIqMvEVAERj+XSRcxs/DLGzaZ5BaXwq91DWOZWL3f+pFZ/lCuIMDGT7ruYkDIUNccoC6MI
FRVEKlfwCeb7vOauzld+Q+s+ZtHV+RVCY33s7heeoL14rz/R2nqVQm5/37GQH4g51jwtkEm7WVut
nYZf/ooMZkhL3y49SwUx3mPMob/w11/sbBpAtbGxf7C0sDg6Oo3yZcq4xvvN62oCS8EMJl5gjMt3
LIMFPgv9w5Lcp4pc4RO9M6rbuWQ+ArOYJKiPAae07lHpUua+oCFG2/HOvhIISi2M+r6tg4H3i6uw
6clPEfJ9aqDq0ZVM+4lHKXgIbaSlV5/kdOni9suQy/jdwTOQGoaFDezjZAnf65o1lbE9QYwk+wuu
bMRzBThyVNckWJBoPfjiJVF9P/SQgWXYxGIpliLkWycoKZWp5f/KocwsOkFy5c3o9Pq9gYG7egzA
lVvh/AZG1ZUuLj1IxN2RY0/CHr3QyQPPpkPo/cDN243PgIDovhT89dnfVrLGA8xfHEiLLTUHHyxi
cLNzIPMVj84Fc5ZnTtHZHiUTaY9WSOEIf23i7hBDu9NiVUu1EQyGCjiKcT/HctL10JJ6hKnndsJO
Law+85mwJREYb2/2XfrvWdsut0bNCLrLEcW0Ste59NHXNf9/SeHxQa7XW91Cy/loYvY5kU6i1ZU+
7hxumXi9lwBQ/Qby4y5lBrKC9l6ucZ1+6tdgsaz+rvT9IXhO0PUikdBMbRoUG8GP3YyrXiTggA0w
TKrZajIBwfB18HaBrSf+EJ8vX3QgnphTvFi+Pl1PnFqNYFn09cIiCXddaHqCmkXJ+Lxu+I6T7KO1
KgjNIml7tGC1CBuMt5/X44jLOfn6v9GbsnkT9oltjkchhc/U6XxcRVKd3fcUC5JyODsNFUIzfj/c
u6s7tFmhxC7k5iTh4RpBBNYjuWAK3yTfWSh/QMNlNXxW52CDVy5JiosA1MR0tdYiJWMiV7yGp5Yw
+WliXHGAvIty/kSB5C5N/0MjUMTQRC+hMIMDnn8TnQUKCkVkKf4csdley0HJ1aVACw3UyIvJxf3T
JC/pOTx9ov/QuGThKYC5ZMKj9Xv3tHDXqvqjWO5wIhr1F3J/jWZQKHQWZD0imAlfurQmRTiUzkoW
t9/ZBzRvncstWO86qpaHUVlfF8rRrB+T7jdHvb5Dd7zWaVp054hWVavGypPXvAb+hKmQyO0gENae
2LhFYzaZli1LAGWNHpC0A6OmXSHv72OpjUXZLTHr+Y1zl5kTns82CqfkpbOQPD70QzPriTo/Jz3P
WisymwpdxMm4/zAkhs4wUcHjQhB7EjpPw9+t3yBhKE0b3L2fbdG2rcnIzrD+7uStvmWQbKe0DDen
r60MSptAthqT2kcOHm++6vnD1J+86bINlvkQ2Hm2o0eOtrvlR6hKUmUCROgNF5r1QY9CKmptR7+q
SX4Wm9JJ4CZD7cKwoys+V194gC7WPth+GmgdHE12AqxYP4nSJUxDPDQw4zQqnljLS412sB3h6c8y
pUueNzC18fmy1CMURleSyIYDrvRow3lWEE7nTGA2gCG7vi15tQVQE1e5qeFx8LfawcrmWl0So+us
6q/RKvW0YYyTSH+p/JoFI3vEqJ2pYQX8qpyAD7XJEFZH9j6mrz1rJOCxfgTFEiqlIhRHcFv0VHYR
I7xYY9tjXrqLdz09C3lswRF/0CAiF9u0/6AWw6HYI9GDTqibM1AJ8jOh71SpvPK1zif/ZayuJ2nD
WCYf6yepChRWUZLJGu5Aa4sLMK88D2qzv0JXHrBAh7/TVGRwW3vGxWgAAe4LLSSCkWN+oKWqKHss
AOHQ3z06P+DiTzSvEf2gmNuevh4taNt70S7fcT8H47XHtVw8WHCbt1oih80HQbNtdD1PJvx8ZSF5
gAzLwkkRNsCOjTEej+6mMOwzfzOtcZw078wm72SnneGRtclFuPpbqx4AXcyUn9Rm/RToXJTJxUDd
q/LMzWhpOB7nGN/nzvjhKiLO3ezT25jwDr4W0YxzVbPyDIzTzjhMCJ8EgHLR1PzE638bjhASABI3
c2me56cbRkCl4F7A/ijjuwMt8BREgugSfxefRqmF1kR5vRcdUL9k/+8pIFOdAMDAj+U6TSSAnavz
pP5aJk4MtYmqtorIUzbddDj0F14FLnlNpqi9r9FHnrga4h/DtPN+coZHZ6wmDquDMHilaxncPrGy
uzkjYlCL1VFFmg8TALnbyHtXSY6QeZkL+SRlkO9+eNqlOp5utcGwU2e5jVAnNRvse6lS04EAEFMA
sJ9/6BCix8PwTz7WOW9ygRiu8LcuMThY+mm8qQnjoagJl5FRDINksIdl/zIN3HCS9XeuTpXpf9zG
8KjITkxESYLHB1aCzyFcEKW1K3/IMiy40tHMbix8sOlToEJxFh0FztogiqwAmgTkzzn0nwGF/KE8
pi8OngBrdAnd1SZnaE4BrczW8N4Rg/5GpgEwGtBXpY7ncBqew8QzEqcKzywHK9MTfUBB8mkumVLn
DwZwf7v0h5bg8gt6FgGdplgKbW/m6AAbb9mLM6NMlNt1AN3JbTSwfDI50s7OWNJf74wAp9Ggu6Vz
N1L1SA+tBPwt4tr0qikkH+AgJYhWd6lMm29aNpBKAUq1Rs/mlWomf9GQB5pia1EXRDYARDI8LyyN
TCMts+fTA5s2xZzpQvPA5/rarS/eQpHTIWhqCXsmapVcn34y3hEs03/UX1vwKkPNDx2KnK7Ldh8V
qsCB8Zuah3oIuPE9E5lshSmg7e/0T1dwsjs7yutgEOONTpMD98+uG15ghvlmTL0miXN8iK3/5qn0
8pU+HkNOid8ZMfGXXGNdyP49di2rvJyD6CVyogV5OQ9M+mNFRKBy87gkQ+k9RU8/QfHyjU2Ih/od
ZLSIMJpGkSAWM8kDEbHX+yY1QJZAWikk+npEaTVqJMT1IDr/hb4yz4Qxmp4b0fYQgGcsRf4/+LJ9
3fbOBWdfn6KzT6KG/j4dhX4b10VO84cMfLuaB73W9QWqms1Nf6zTfcBNxH4KWnvfI9TzOZLiEGl3
f9MS69SJdhrjDnl3+y4RfEDjxb42Qr8uUr/zSLca8XY+vEyiGcWZTgIRqEvsHNMzLsIhgYWpaXgN
GFslU4HHmTEwogd4ioaux6TxTajFul5KQ7r/XB/BkIHK+riaCv7UQW0TmEngBr3zzMOfIr0Adh8n
EkO4B50GDawnCWMHae0fPSGbRn5Z1/P+1i+LCJYueHHou7A7Fx9zhG6BlX0yxcurSqjAjJWk72Z6
vgU2JJlZ4Yg7IToRniVEnQLHzotg7h0+wvLTTkZ7vLy08UEr4qhlCudoqpK8dhG75m6ZGYwJZfWV
DfJra/uq9yt2vAA/MtKuhCRI7ZZ2k9UT+/jqAB7TUkRjjk+MFbcBI2BpXd8LMSBTyxJJvrA9DmWA
vr2H+Zgym/6xmZAKu04KwZRgEfO7p3/RpuMxoATalSHHZPTrNal4smFLu6EnUDEwO2fOwgjcbzwA
r7IRQun5dBX5cbd+7WI5nNs8br5eg90dLqcCCDqGHAA9KZpgMIBlS7+AMLge7DNn5lV0jiuUWKHR
/IxMcJnIsYMntcTqGaVrVIZp3owbqrZQUY4Vwni0ueF8k7xkExbmp/ALesOOd/awtGXQR+RJMSkH
rpkMxvf4pOjiU4esixWTTjghe6cEbocEg0L2C+KKUBec/MkmyzuuPh8z0OfXqDgfl+2Ia07PY+rk
t6K4S7P0F2ni1HTgCMKopT7P9E1X+IPV3uTYcYuy/dfBnId1VRX7zSmwH94ckUUJDeth+2fjRRmQ
zpN9NaoGExaNIi58n7KsMJY3K54a3fjO6wmsb/9ND9wRigwW18FW3gBy8ND6zW1y0gtcvektLXjr
au8DqWzrMSTWTfZ0wk8H5MnqTOQLyjEmwwkYQ2oyDWtlRAjmP/BOKJ53c58uqQF7C1isxJikzY9D
M9gBMuWgqWGRhLIFcd/Bm5tv/kdCUsCSDS2j+xthUj1oCX1OFAmv96KLUHurNr5MnKIPy+L4asEs
JBePzdI+G7qbcPqkoyyf+bvgjDYWVss6LKjXDoyGpkxJlMTKyxMtEq3g8JRp3P9YXdgJBxY4S/Y/
YYVibRkuafE5Tm63AxyZjQiZefN+6f7Il9VfWLHsmA/Pq8A0RVeP8MCF7tGliAd+eB9sNHgP6pPa
DXFNdZC2ma4V1UvrUTpzmhmC1/Ufr60b4KDJr9uTFM4tvc2gKAFl6h/DpgR/JCxoYhaF6WwBEvAE
iDport4qMICa45eAg09MmuOenIN1XK1kpGiCD0ly3JrnmiUdBb+KAUZEcey8T3/QRX5FtCl3RTCI
Wdx2+hqD4y2pxZyk62awyHlrjBYQARr2y8drNidPUd2CqDftcKmm6l/syj/P6wsH5udKgq964oxE
tFCqm73rftkI8iykJilCC3YXRyvv7okAuy4NshYHH/qNLVc5uGBPMvmDxYLkXs/9ghwiuiSiSel3
Y/jniXzCDOP5sIwdH2UtZbCn1k5c1Xo+O0wHKu1EqywnPLX/S5AjVZJARBXL++J4V2B5fFYmiBFP
8RGNtHDLWMcq6uap/4Yx2nKnDNU0rFSNm5bHvHonmbdTbQN6TbSOnK9drVsLlJqcdvHUZmyY/OI2
KWDi7VC5CV+BWg9vHMMK3h7jhmaZRWRRRJ7fP42i35zvx2AzpjjrMHaYjeY8WWyN4ETLRIl7yMSu
/I4EAIegygvKQsDqoj6bHrxn1LvN1iTCKRhDYtY1zzilPuoZhvCRNzz6kdKuVYJ+mbyCLfJbIxsT
9GX9H0yUZzIr4itPcexKKiiCSwwIxDBrr1COjbxb49YzVF0ovIG1TBJISQI9stZNRJ6DcDuCwo2T
Hh9i7xVsEGGTf3dcR7GAPpZDJbS/9eBoP7THB0eg4f57yewm5FBpFcZ5hyuY3vp+X1ZQBGBJOIKx
UrAj89tvLOpCJAhR9uXTErGjqKs1S1UKmcZIMqlC0mtiPwMCm485wwBMOx0+XEvI6Oo8lDc3Qqds
6AHnsLiKTw06/sNNBZo5IxII7s2pPNIkTg08bisIcigz/p4BnPuNkE/SEDCRVuF356PJD+vxK+Ww
0YPie233f/VbeF19/uxZkNPoNjDTkg+cPXncBjk01at0KFCpyByibgDJBxBJpFjZV4M/uvVK3mEh
cbIfIG5dDcdBKz00jO2aOYOw9LTFVUoygOBbX6IEAclNDNJ/cDv5QyxVDyQvCxjNYMwyi3N/Y+5i
RwsfQHO9RgnsRpUE3gkJ18tdQ+2KYu0E12AqN6XWyZ28iaqFHcEzmXHPjV6WAooQS3JJXcW/umRP
JV1GGOa5jGUozdWenpdk7EsKOA18LzrFzLui0aVRisRscsEoVcu9LLbygn2P8xLkpel8G/7Er4pW
3fOYZMIN34pvdYKPzeWZeXbsEprZCOQAinJT5lSBPnCyOKbcjKs7TyfqQef9xGn49B245BjCWXIt
UptA90h14TOFS28nSzvfQttfuaN0Lq0mcDk1GNYye2SXGMzZD6jjqa8RTx+oilCaZWa2zlAJhUnw
D0Df+KVWoAWT6/ZIkL81q/pppm1/kG9qTVInDxzliIWy2cD+lNsJHnTAn2Zma8AooJpOeKTNffxw
oGy0psFQvQ5XRX+aytMeAbIhZ5H7rZuwBR/jvxDZj/DnCZRLRzUwNrNVGPJ8HVTzaa2OEDJshwHF
sdrtx7gQ8dwjC0eSIfi8WgKnFNpP4U8fe3hksNjVI4CzCt8HUjozluwHVc2KdPynaS61BUEjyOZF
U1pSlLITKtEm3DPnLoOaGPF0iuCyuFwmMCOQrHDXcqMFD/TU9lcUf8rGB6Z8MNVx7exdVIw6rPGJ
Pt0kmQMQTXbVhMxecJMey7l1/WSltFmL5z+5DDPNf/MeV79dELo5P/AZfAbZ4nQW7hop5vUUQhpR
VMIkP4oiC4WizZL5wJhXamNXPTQmbn4KBQguCqZBBV15SoMib1RkLGveao3tYWdXfr/8TGxjmmiD
1CvaULhuaJ+dGRg6yWyOpUDrPxK1iNjxqKSz+0npad08yWE3YgARwjkNn6ijJr2c7FO1l7weZlgB
sC5euV+fAf5+5LKxkCqBlTf/xn7HAmSiHWdUQi8QPRIGXI1sjeu6EYxBVpVgqnBAWwJ7XinWSbl0
25sjY9QJHs046OVxDzowAx2XvugkL+EjuZzsJPnZcoJUezzxsvq1ZNN83hVV+D49PH0PKxxWL+Pa
8l4HHF3VtbDqAgyYsdwF7s60DGvAXotDV2y6tJGy033hk/GRlqhpbFs8rKgfGGFTb3k+BEiU/4R1
rr1VwANmDX/5+DmIwYj7zOM785XvXOI/tsc58XEHRCt1NoHl1MoiQaVNY3g3YdGrTxoaHJzbPvuq
QBUqn1K21WNU9SSsaSrA25PSmxzV8W1SPlVveudBVIthS0pOVMnoavVxItgduAWB9+sm+7SsumXd
uXkpa5/tSEdGxB3T5xQfdycl1xjYX0+xkGTiyxPHVPsxqZTm/qC6UrB3QWcGddtTHJ3khy0130h4
v0fodba0zPSm4TZFCAZ+QjY9jgUd156LgPfU1Sm+im47FZNBpNHRzsAOjubA3dNKyv2/Xahh+/CU
livy8iWmdTKqTFTf2cHZSETlPTSW+5uuE/XEOYDC7kwddnNtzM1FQY/F97wOo7ZWL2YWVDAHhrnJ
df//Uslr5Sx5tFB7sEO4IygC6IZAF/Nxf1W5FeHVXiNLQh6DU8mRi6L8JAXonhEsuu/4xH4U4P8i
QikG415oCte/waCoBZgD7HfGKi4mdMN8JbY7Kgrs1rNhphvE8753bpCZBmnNeOCkGdE3aQu4Ghfu
YvYbWQVtH9QWdaTArEi3FwrSVCMWN0gfKsjTmh/w9G3YEOez263fhPdWboBeMPBztlkdm6vI/x37
i8FTifH59FnHjg/xkhXHO7lDQGCnRTrstY1wosghWdpJrWQw4e2i0QRSdtBFwwjtwu5poNAlswp2
Wq4OsKcETOo+wDIhOHaIOq3ouMfsyLZ1DR76lRqdckbipO+PfOB5PFxJYE3HIgFhlxA6xRrsxKan
fUjScCt+bMOQWeuUehE3cfCNM4eLEezGL/KbDzRPyQoeLFMUUQk/0tZp/Yv46nz0IDwKVlJrbKp+
JrIwT1iqLSB1hYahRodXYQhXuppz+xOGpB9L2eQyn5vem24v/KlU8Q+bn4LPyekfUBE/oXOc3FB5
i92cKuxvQ+qjQutCU3aUS0opFSB8gF3Prpn4nbUhZ0d69cF1pNHpJLjBbUid5swuE+Kgh2plL4b0
XgrgOZ7ZmrYS7ouJidS5UH/D1DMVvIN42cflMJTGrfHJG8dgUT5TJsL1oTVVXQXB9o6ye1GOKbpl
BXiZA6n+YWv90fqMe+/fsu4WoQcCoHI47/BJxmT8YQ6gx+pKSSkVQ4AqHSw/O4dyaXJI4VDbmq8p
monD8VEVAcspRn0RyEV+eg7LZaJOaDQFZZdAKg7nFN0imF7jiytSU2xmHOYfEiHJASVJy+rzHLlK
Q7/FvzAWhBWR84qyLWQL0GBQqJBenX0GiDI/mGpvBrwgdu0xQpuTqs0HKGxtMLiDZutKDEvw2mP1
8I8makA6txorXchtWZD+tgIHmCZz4oHA4QMSWyuLtVmjTnomHweDzTfPH3sO8WQwY7KUko8KUowi
Yc9V00prWqeHFyTtMtqnxTqKuCh9JCIUEJ27kS+j96IxkHAu4MGBbS9PQro3IwRaaTyKs3cUaAg2
6HJt/lZZAkuA1lyVTZjg+jwozNkUf4B7JdsoNNRuf7N30G2zFsii8Cq6xPLCEQvO9Pe9skFMCtx4
370cIKs7LVpICFJxOHCAyVNk6XBGR3QlTk4zBpAePHNrT0E0iuMrs7mGeh/Y6Cbmgv/wy4sYLypk
5OZsSQhTmV1UYH5SyG/zZbHI6ysgsXzeCM365q9r7wcqnNRfQz7nJlE88MYSwiNMk6l5ZYG2vwQJ
8UzTrkVikRO7PsGaX1GeaUqRfPO6Zw6CSWcghOsajdNQ6H0Bgk+AUWpYFazkl4tLWPXZWXhkxX8U
q/elqU56HAumoWRy0zLy2XdJskhZcveaFePhy95gEnl6ONZ3zfzXoQyM3E3/h6sarMyb1amYnN6O
656TjsOMzgZ7t5AQKykh5Zpw+CYhhgTaTCEfJMroWLkc55sLeA+hlddU+feMdXRuEaHkvQu3HH7Q
fxXMv2PeWH2NhowXTZub2qLysZyiH3UeuDgY23MxCY42WCRfkN3PQR5eYPO0BTDQYB6PNYKRNN2W
4gCAbX85KDLIFdz7yVQAtQJgWHT5WDTZQZWiBheovKqKxrVfeuVYG3p0QS7dRdSua02T6V2kPOca
nuxC3Y/a30Uv+uX/sTnW3smmZsxcCxJbEmu2XqQIyNhXbFlVEHJNP7ZqPmaXb38wqi3ZxEjTjSUr
aH1WTdz8jfKsTqr1K9vwokXeIHd0d6nVbOoK7UM7syXbKaQPktQkqpTuSSthGkDKQyla8EPsR59d
szPXoMa+Tgm+wgPC2yEdzHsZa320OMk8UW5JAWIfN9JU6YMNlD14EH1igKh5fwIGAZ/vCFOWmw4X
f+vzcEE/TgIMoT1F2kOcQWNx9TTQ5d8XDEctgFRLpnwaU3cH6Cu0JjkHiecg2j81gyfIGtP4LXRd
qvu7DCanx8ZMXdJWQhTpwqARGIzuBGLl0jGVZVgJfD4VmAeePEuaz4S9dv46V69gYtZUTTAOoxNJ
0MD0FdHaFUt4hpikL850s/1FW/y+6SdmuK5khW7zQaPA//agaJ90incbjwmMq0227/c4il2MHmZW
uf+2itTjN2KG+g2nrSeM4S5Q24tkUlkBdnQR8ngZ+YnRLy9VPTvg2eTNGs/I8SlSJQy0YxTjgTFA
gYK/dXtvEpkGGCuQkKR6FO6sh/2jNdUPRYLwjyerKHhNHtSzTm9ug9iVKeoq5KYmYRLGYHAh7Eed
D213cU+tuwT/MBVq1VwxVpk8v2DGrPNYBfyB7es6HL56OVCNJ8b2Qe0ZDvLJ7EDNgnll4TRUDzJ9
iHSiy4HvvG1oWrxPpnw1YQbep8OxtpPgl/QONS4Hn0pyDIO7GeIk6eDGh1bRj3xfxxIg4mSZ+Tpt
m/2Qc9NliwXz6d+cFmpBVgOZwm2YT0z6eCXSQc7eiXAHExQ77uqGCf4wrHaXg9nSpxK9TrKUIVj5
roUE2t4R25PnI28GX762fRsT1D/JmV4p5vs8FSMBeJzSyqv9h1rrmxLafKpcAcnXvc3dIynTYMzU
uDjGCI2q0Fvkb0RTWlAoFoa6BQvdT/P8UMXx1aE59aVw/BouGaiXVgUz+rlZhKt3TTmXORYDED/L
jYx2K9XTTyv0D91j0v+9nnpqrdhs5rNdcjeVlI6dAXKMzpyz25QWNUk9LhJLM8GeKcLQMIlyiECi
mOTIX/h76y4urVMrHck7SoKuCQHDi4PLmGtbprpv19QfjD5gU1rtJ04Q1b55x/oX7WnI3Za+phON
hHfysQOCXg2TTbV+r25OE9gHX8KhC03CH3wOskvi1KDJRaintzOJVG5LGk2JpRpev5X6IC+Hhwl1
kCiHT9+4msgbRoxdGzSVXQJnNbC0XQyy+I6FMzHA+kiUbhKssS0dCyh0QsQxlQBc+2OXhNeWYnTP
J5IkXhUBlFjZXeDDS9ZZ2WXNkejCu0WkFo04q/oCBG3pHUNu8FuCO9dNlEs5StKVEPEF+DUPKUZC
Mua+Ur+4AcUh2NeN4dPKy/oLkY5bOIz+xio/e2BvHIBoCqnfFNROSq5KDDXksQXKSg4R8EyI4qpI
rKaMCKzMqoDeJ4THBi6frzt7MqR5m6olFp8Goz+PphWF0IHkNAoWkOl72eXcEeyERsQ51L04U7dr
IypEc8P428K7/IMpfuC1bicVEFCrlFOsaFm3kBFy2eSeeRpQUER1yELSxluTGClpMB7KYIykbQ5y
p2oNxsTTbOTWH3go0phltMZoWcZORhF8FPG8Y7T7vfFEld9sMN5QuSsZN0ug7taUAT/vbF4RvO0u
GCmDWPJLNLdG/CwCXoV23U8WVpNIzubwyQrhKK6QO6kR0KdqypKxfLdF4G76Q/IQjPCLwYGp9t1v
UmHFcDkyD1W1NJFA/Y1RWBnlizeKznGYj1D4t4Q/SD+Thil4Q8W32Bka1ftSOAo29+Om0WCVJEVx
ibSTttUdIB5YFv4dx5xdD/Kyafd4n+klOKL1mu9gwoVxvGeT4VW5JzOWAXJX7ngbcBFqO5fO60dr
E82AYz0j6kqA3r1MTl/3ZX4QKE1hKqBWfkYgnAscQkyuaxHV+h+ij6KbAratIG6LhPfLP1wTRZFn
usykTS9KhXu/i1gvOgwuE/I+9ZE/Bz0ugd4t9NpNbv5yRsua5G4MZYcrYP4agZAV9KbYmbV9eRtH
pzM2W0uKB9nn8jYstsSSC2m9SADyBDEmvLl/BNQJdhi16bF2+7QbqkWnTsG/Qek4Oy1mvqfmeTzR
enfyW+JoZey0GXTq9dLw34Uhq+y7+F4sD953sQ4+lujxfK8rldSEMt61JEWFc40ctj8ELOw6lKBn
TZY5n7ZxyGVC2YTKuXUiJcZEG/Gs6QdWVmOZvHdknRb0b9mHSwXlF1PZmnAMQ1L8XgkAWDgBz7AI
s7D/i5UQ3V0Hb99TO8Y12O1VKslf9sXB3C6qLY6bRj8BF1CNjmwRZpl6ZNo+HL4o/4ATczjMcdWp
2bl3xqpvb5evrPiquxhWcM7tQ0ieHlauiVsoOSGnJHn+shopCvxHf3084mKyJy5jWWN2Irk+6boe
4kmkmJRrhmGxLAngEWw7YG614gG//qY1l3EOv+3DJYrraKHVdU/Q+InMej67TQ4WZWnmb6amx3X2
/8kNuN427NiO3wddPjCnWw1HZX8u4gBiffGYkXxX3j/19h2vjIp4n1YXyT8dB+EWlCNrEXwAEv8S
vRHmMzzDwbwBeEiJAS9yflYtCWdeqBE6O/Ph2BMjbecJabMdPTdxiaJo5EjTnJQJD2oc1cjGpmus
0gDie3WVHyF2nBD5uMmAKpojktq4NrTqX/W0D4EnmCxQ8L2JDYxKdeOPZsS71auiyPBVA9ASsxy7
zWKULxGwQ5BlAdVOyFG0rXASqgDqPOWDF67bx+ThKtdPAwhbw5ZunjUp0bUjUEK1Fa+Qfx3e2xLe
pJwkeL9CyMZGnLg/TgwkzYB3WxOYQUcBZ/HBwINVY3uR+vDBR/RIeFokInwsqAxh/aVAhEKaN0QH
kPNjBfOvuywuLgpBoGuRcFRTTa6ifxprdKE2uBLuyodUfq1naWeCLNAAixJNA6rTyuqSHEQ9GsG0
A/sT2qlH1XeqC6IkxRoRSaiODuRF62c+ehTuk6Uh05jC4+3JHBg2pjiUpI1nDtQ//m15tmLPqxF1
Cs2c4pNGgrzsthe/hLf4YdXURA8gYoaqaUELbcmGnIUxBSrlVxb4paoe5i1JnAHoMbtp62PMoJWw
4J8hBC5YVQ+gqLfxUR1OhVIl7+75Pkn5Csdc6ReFUIeYG54aDMeRuOJKMFuPmn963t2WAbw8CHXs
6Rbd8SsnNbFEqadMk/RdfbenKgeXAZ2oEg+qAhPfyrDmDtMw5Snrlqw9N1q7rgCzw0Ge6cmqrnho
YDJklj5tPEcGaI28QTpV9JlcRgrpDLJxNjdcICOmvx97dYlRAyPiUV/JwVLkNcwOxJWM018FanKW
1ClVBW6952ZT3Nh+VzccA8qDVizLL86MxFltjO6pYbFZFrZk6gkC+PilLeyuwgD2ctew7D98KPNP
hDlKPH2Cdo6UL38h+48F+SlmRQ28jVhkNEmgKK7IF/8XadyKYQ/t4juPCXUsqP589swRYD0eZdVj
ZFErTZYNMDxib6ZeBqJU/wno7z40lyEyMgsk/oLgGePNihhX2cnvQTjM7O0rkvy7aWjcHnk61JgU
rHGggXl8ZSnh30qehdkqxKr4RgNelHnZWU/gHgNZCQyTvGQgtKL795r9CUI8Ci04nUc01Ds7mceo
07GjQPqEscA1adbJX/SSPqleTVikYgfcb8mhGtHM7N6u7AB3t2xuPjgv13+AG2eqqXUURiivqJFp
s1vUHOFUmtHn/tGyGAnCFQgBFIZNsT+VHZbQtxvisX04I5YdNwJGKLN7duuoxi4IJAr43QDunVPO
TR0TuHyGkAc9ISlO1eh4phejf91NaKQFgc8etYNnEcFct7RSv9+6jV80obO6ick31Pl4OPJraktr
8NA50vdHdBEL//3WTEYulIy8panLmLnguCu9aNMX/hOG1j9M0AOJ5XE/2WUW0ZDrMNU7NsdzD2Oq
SJhg1x4M8Bs6NGMDuMaG38Wl3zx3JlM7xNyk1Gc+3idwzGuETwBPct3u/s2HQ/4tB6DDwu5UcBUQ
4DPNIRUIqV6EI1ljR7SuvaGCHphw+gO2RN35alEGcNkCJ9AO5Bd1isp4paFraM3G3unEPJz8il7M
C1Yw5yn7ML/tiuSx5rC7Kbo5ZURHvK64zn+aSgZd/2sUiePWJihU+zvoPb1MSHySdPi32fr6eMS8
dVt1EFhsoU437IpBVbLPikbvro9azdxprX+jQIeyJ3EIk3gNCxQ7J3AL6FelHAg3BQlyfbpHDol2
MHwQusCoWQjmywKZdmLuPSSBrzgPUV7xKIqGl8duIOwucZPiPflhuZ9zJkiD2Fn5sEvEZvhuOy7K
CdGVNsKogVz0cz6GkypnLPS3zr7bXTmzRPo7Y1ON9iPXIjRo0E6j2KajH7slo+u4lbaL5X+Neyps
Se+V89kuWU/KeWZkVrfMhRDqV7/vorTbe/txHaP4oDAabj04UpF3e547O0c6guc+Q/bUWi1iewyA
cwktse9UznBAhbsBF+Vu0uZEtXV2sbtzbrbbO15mLDF98moeirT4tELTRRti/052/nyJsFZkPlYf
eD9FbBziPlogIykZg613kL0RklRmAzICrapg19c+k6vHsFiIDas/6a+Pla5VtMJanyOsTPHoos8b
oYTyHGbrzsdsR02iTB+MzkNmL2ng62MbfGVRTo35apQ9hYjHthtYKDgRHTLBJRJWcmQowAWrF1WW
AZl67hUIXtDqDo4XQwnTHTUPF2lb2FR9itWDzvWbCXMXNI7iS/s3Wy6mwwI6IRzOPBw+CSysnJQK
VDSQsJft0tFnwXerpsnKt1mGfxkJJT2dSYxYYEdheGxq2hHF5FVtXH2PSPtOwK9fj7nRkiLbpVm+
VsgcQP+yWKWGpdcQJ/pdwLiX4rlv0EycVys79Oc+uRMagYhXPmdNysumUpuRlcaFl3ufDy5EOZ1A
lYnR7Oh0+A1FngjL7xqTwNXwBvHNaZnQUYzoU4s/gbykJkrKnuSbPqJE2/QLQZ8/KLogxnhC/KfY
ncjkrJSm3/LfIYfafeyqY0z2grvxquPB8pnRfxzMeGm1nb1tptnekXZ4i+nWE/LwRCu6SAsnHyAw
pzj0xUfZs4Jt9eMjg1LO7E6ficVgLQRtfE/1ltzmt6dc9YO01V1BOCpquu44ZKm9OdRsN+7PLnDR
Jzdz+elfQ/KIuhdBrZgkZ6pctNwOY9OqMMJMtpl4tKdFRAKq3Qh7uLEede4/5WE7mCYWK9JijoKJ
xVUy9ZhEmxGhQe9w8TU7Fr/QU4rZh9gJu+ZuNmq4jAeZYtUeeqyjlKE5vrfWkybBz1PDghRBFmpk
9zHac6Ss1JZ85ihTs4PA3mQRWHnTeWQmJteidPNKD8D7KipvOLeMNu7f8h4dhZOoltITpAjaB6JS
URTNB4j27tHYrc3U0WYQ7HJEm4UelA7T/cCV93Z6xnVHUobFr7x/zJkTN2OGEOhojPAdOPY651Fr
j+LxH+VCXju3kwuXEXktIi95QSu/UGmOTIPhkCBNuiAkg6EUc2Zx5bCNsrTdIjy+qKT6kdtqg9I8
zBozMcLxNpUAo6qvFMK4uIxJ2PhIGNvSwLA4HQ1OAX0V4obbvEdUL5CNYptrrPGLQfOUmwj8utzP
F0wj1pvVG99PeoV5FRRX8jE6ixCti9wOq+s4uW+59Q3eO1d/0Vj/4/ztimPGyQgsKNUbem41FWy+
EaWlvUd1fcz+v6vu8gbRmE6d9ACOGebg4kxVqFw2aqoShM4Sql3vtZjbmYCkvLckiZvn3KRhKzUv
jZa+iKcCliuvVZ+R8siu31IP3v1pJQV9PVayB+z3YI8oVsYlaeBiTsuPg3sI4krd4edygQVNP9mb
7wKH+oN/uv9ZEt4XSH4KxtJstE3TFsDaLY2fUHxX58teuM5oqL9rlsiJlcWuc0TMu5XsAdCo2vpw
wfJaRmdxWZqgPx6zJXFE17E1YVKhHqV/8y9hy6KABRDLhsRaCWAYABSaBuwbxx0za6wjWt82ztVK
T4b1x6nX1a4/3sxdXZrmyI5TpdPrTFKlu+b5PwHrXo2ieSpVYgchD9FZsD8hUL1HmmukX6yAnopS
LI+ejLMVFhwd3pMzl937Y4jk03RJ3nLqNWr55dHYblCpsRA+JIeSE7mIrKtPS54RfpZkQWlZFJhZ
QvUThA7AjH6D7iD0ehKyOhB/5kTV+QRnwrpJtuWwf677+5MohxaeGTZb6kroPj+EyrqNoIxogk1U
h0EF3VbBh+8FCtIL6Yazr5wV5Y1ITKO3r8i/VTC+aqSeCZaW/BYF09BZ5PgbAUOtkqpfwYQHS42T
nhs2po7yb9jTduBE2lybjxyr0RlKetxOv6ZUMtRhVvdxdtBCFYZN3KwFjQoWG1/9dgjJcKcw8SGh
fgFtf3HqOzv2teJqi/w1RxzQW927VCmrkdl8ezKqmqX9fT4ICnlA6wIdlUwO7jZKVDkL17qRMWHn
xa/3tsL6kx1iAeYyBhB2fMJQh8qbQ9hZeXCV8DnBwvbGIa/1Pa9FASPTYyHfDNW2hfH43Fer+qor
v32FOfqcaPdKqK65MuSacSQpq3xZxHdB3E5lTtvnJo0ehx1YJk7/cT/F0KNUhMgfhBpXO/c5pzG9
DNgFhfB3PqX8g1mDiLecTOPNzFL7/5CJDy3q5Tu5yNK077ILL6Tpv9SfvQY0meVPC3ZxTpsJhgHW
gXLSOkN7Fw2ZQhUG8HlV34VTj69XEdZuiWa/8PaykWpEhwozIrq21bhgto6a2DxlB9Jo8YKlNPK9
8iPPk1dvK7FBh57sRKfwAMUwWHycKgTQaA1ZR9ltjAWgGwgrR62T4lfakS3MeHinmxozQGNmbtcM
Q7gIdkd0vZix8Zs43Ti3fmeboC2J9i/xvdREvMpQ2P57edt/74oO8NIp0Sr6hG+CnE2GAMjN/2ox
Rcy/h80lSZEuGiwcv24g2SmlvnJJsR3CCY6KROA1FgUKKswnwK0Dr8xFbjTKxhlQ/pM5IgIchUww
FtMgs2eyEXKC6wFeShw8E0XhhtbtUDYkKCpbECzFNlz7b0Is4pzwRc+rtpdrj32Fa7eKCj8p//hK
Bs4i9XV7nI28tjccLkaBVxyjfJEtv2fyysAVwmb3JzrTN1xkUfqLX2tDOfr/dohYU1/3UPnUNmVn
dM3Vj5qNwcLEabwKtXLV3kIc0TQvpULpUkI7OoZWR49A+yNPNmlPDSWcgMC+Ffj+Gr8kEAYG9Rkl
5ac5glfq/KJZ8GJDHYleTRZR1mql24VycZaVXGtG22GeAC5NN+LL0+4ZumFNFd0syxijB2aIHi00
rGZkSEGELpWdjnmkZloU0P+9y2V2BQPBIVDZqFE92oIRGLSLL5POGgUR/6ll2VV4HuodqHn0WKRF
cD6kCcj5d7cfddaovYYXPtn7k1THYv05EyUb6wRA7dytj4perm7Mt9sd75ieGjneAGclx+tD4PYG
JGVw7lFHibm04hLt3pWmdzrSwyWjdUlgl4NW6fQ0aLIxai/05rp/fIjehgu89W7TZbrcGs4bULuB
Z7Q8z7GZUknasZ2gUD6q8MwjiSlTD+Lw9d2ChgrDFKqvQiqql+dpSmv7zzc8SCzsPC1TIX3Q4OW1
I3a+V3twHUsTWFYgtD5VP6iQ9Pgjix9fTEAApbQRHwhEOfKCic1mfwl9OIF5D1LF5iwhhaRC2FBZ
33O10q/yzIhUmQfS4ecXXOFb5Tjo5knhFwE0v7qEcQrUjrf1Dq0AqLq8h0JF93As2785yiMFBzx3
hN6j2zF/nL8j53GZ9BXWUZAeW/C1e1DwAFEe+gorbg0SIWae/2AKKDjis/4wbT9SG8RL8oPbgBHb
gJamKaC3UtQ8mD75avVgLcJzMGtTYwjx5Stmyox/eZw6SgYuZu54J8S2brWulaNnB7fvatCBWKzC
KqF+y7U9RS19R9d6eaW66N7ghACqZRSdN3S5zX/pBh8t9qewfCDJigSTdH2/2mCHythPsupKh0Fz
x5zifVRqgT8p4a2kbvTESweflNdZSqp6+/zGjXq4fXfv6dA2Lf/BvFu/HxyGqOOcTg8Ug/y+DGPc
YqGWIWtSAQR3s6Sh5ZKsigYK1DxWiP9g6v23pEn/sR4u2HYB0OxJ0xscFJa0FoNSIqzTNooiPSnD
awr5y9Sh3jzlAuIN3RzdimjyuYzif2Bfnnv3ltpiZJOa5SOA9bNJm0eQp92XPPioFUF38YZgrkIA
m84+P0DfjunKve9+pww7ttnsMpZpk6B0WfuIvrxu0iRlPcljWgkyXdm36GF6gzqC0xqS1PjG+Q9l
NZTpjBTGlaAphzFJ15Lu0bgYeaUZTK52VHaqb4upt6YYosnpv0wbheFl+8ytsz+iP1j692F/n9tA
W0bV84/1K3o1HcSOOQsQ5wei0kybmM1ZOdHU0sH9jmVw4ohcThWNGRvNkCkTZyhZkPJK7rlE3YCR
AvS6h8oes2zjhQBhL1AK4dX9IkcaASo+pTVl2slWk684r67vElZxavyoeKlOsp4xBcNdzoEgRBPo
PzZcUcNIHffyM4oMJTpgXrav9ALOw683EHt/0znxEp9R87KiW4P1O15GyFbSPgkD3cfXeU8Gq2TF
Ps7EDWSl5kedtuZb2BB+lszNKn2fiPBpI652aCQ0a0+oaYV8Fc2kOZeWy16fYZgTXIICnE3MURa/
UjyTwZwXsOO/G4eBzU56m5O9nKjTLto1NETrST4wDWG5kkClbL8D4c2fD28Ed3jIBkbSMTyu8Iwj
YkSfEaRVLzaBxCT+EAc+LZtNLUJyT737qDyOePBnzIeBIq4qWfSBZxQbnzmQGKPTt2J24FW7Htmq
DvtolX4ZV6jx7uHnQ/Q2nL+q2Jq+8cPws3viSGW0EyJHN9q452khd8I/2kbkjbi+k8e8JQr5Ts/0
W1pkXIp8PEkmHHhgYQW/6ztM4J7JcXNXG8DARk1NEYFmDaQcXDSFhjWmW6b92MHK2ht0RcApBbzT
TLxdH4ouwFsdrcmCB2ut24dwH+OHxMSHb2FoiIZ7FwkWS66LBeTYHpya7MLoc9cTNPm5Xt1pa9qt
//BPSDxlZIIRdD3+kfzHOygruNRCIfDWeBHULandw0cbCgvfpckQEsRxKN5Cui67uLWhcWABjz5S
QQTvPlO5tVLiFS5gZ18c4WWiN191fNofF89fCfnDSdYCca9x3NTcPz9acsG5arKYfMAtTTYes7AT
NhSZo9GPu/AJXV0HIPqBW345ALv4rJ485AYYElTr+nGRByO4ZFo0xMTKTHabYBnsCyPQpmzPTfOm
W4ayw12mXR4l9FZe7bktZfbpd5oSdh09O4Kh4wVrMbdRPh2cTg4xqBNQR74yu1APjHh/DxWH6wM4
lBTOcV9Xetkr0iXwcFL3fcQSdHAbzYBPmAxC56u1OhCiHDzKvshKbvFvUfkv2AmI88gTr1EsOIV4
RqWntWX5bcnIlYOuXYNNu2wWT0C5uUAFCwAoo+D2u0YllpGX6gVfUz0kx2Pq0YbihYJD5JY7OxRj
4zfCVy8sEKoUYTMVsnn6OxdbNXVUJMDwkKHl06t1wN7vciXpmmTOfjAL2U7OlXU6sB4YtvH6CkqC
xYPn8s43cR8M7Un3qY131rcKkmqeVSAgwIo/6EwV60fgEhDmdj2UcM3w6bjW/6EeDvXm3N4jcP13
SCSMHjIx+mWBg5skiyBDFLGOlQggd4b1yCzuJaaEOeRKYqoyOH3UYDH8tfuCiPOo9BZnCszugYrm
ZYggHgYib8tJ/peNhJYbRqmOFV6x0DRVP/VAb3GSGrCg5k5u4lKWI+sJc2J/IHXnVpF4aEE3BeO0
cE8hwDxv1qlihNgg2BCkNSy+MYBbDH555ER3VDmB2NPuy1SR2gHP5vJ6Tl/mUbnqJcO2cai76fsC
uts9J4FJqXoPgT7WJiO2AUgjlPDjl3NtPNq/pKAuuD2TpAh7/kQX8gHMJ3lk+TOeULjKS8wPls+N
RszpJKWb2yzp/6OTm3EPm89dit1/+UkM9690RajdlUfx3iJRPbKnOUwH88d7qRLWmoAi5DTfUXni
QBuPhhfFidt76+DkiBL0a+uMr8WpGk+M+mZ8MOF3C0bFjb2hJ/OlvPp8piM0N+nopVBvvrn7kFrG
QXFCF4F9YLgRjh4D+t2jAL1xPe/kLUfOmr+GQ53nu9VLEcoMoA1rCUSmZ8ZUx2+G/T90HDagLBln
qli4zwQ+jYKeQcoPePgGK5NrAM41Drqwe1cb3q8l9BIB2GsphzqrdfZj5Suz4pHGCrvPRH3Vbcm1
P9s0ki+Df+6td/1vPLV1akj/n5Igul6/luFjEAwXW617PZ08ehIZGPPo6A3ncd9KKUeo19fdEnHg
qu0fCpOnboqzdVTn3IUMkhZ4UX90VsSCcuFi/KwyfvlkJX5qHNI8bR/BdhBf9HwdYrlDMkuK1DIa
XrWbkFpIAhIDGJuB5AR4GRadD39rB6SGsYiKJ+PPNInWtKL6uNNj2Wb/N0UVwtzskzjdXNb+9PHb
OJBz/oBVvOegyPgi/+BRmiGbcATowMujMWn/U4FYT3warsCuweQw/L/GCDhcoXOvYA0xCWwKlgyE
SVO9jg+cvSVszIKD8dD2T2jS2QmXY2AvmZnd766bHkZrzrI4oPxRTW2JHzeER979N/C7cJzACFQw
Yw7VS6FfAJbvC8zE/WR1h8rr8nyi9RF/iy2Y/XSqPLcQ0qFjbWY3EzLOGhmG3ItASJ5Vh+RQdohZ
EaAGHDpRII0ZOyzj5HyAWdL+wNyGg1O/Eg845r6GlYUT2XqlSFCqg1Db6uks0aCXruJGjDGPKAel
CquqQjZ/+hlUfWCHxY3Q6IJursKgdVYQljJdLig73f7P4s46z4HeTnd3IoXBJaS3jiTJXY/potD4
cFF5c7dykM3y7Bhex75o59jlrUNi2eeCLjB3smKb87qg8JjOYxS1vglaPFanIEtduPAbP/kb45OX
dc3nHoLaGEG16wydxXepuk+JgmZFcfezQIfn6Lo34rN0sUsrGVnZ+88hNLvkiZJa5FX0U7yC66TY
/ArDbfC50q4OYClqDBmDJ1nc4EdyZXKTTwZEHcC1IlDK7ZA4AHf/+c87fSfTpiA3OeAzkXLAP1qD
BY5LT18oiTeOYxAmqGpHPe0ghbEe0Sj3ouR/KR7uiNb558KrqziEkh49wNQiGavWOyf3vQdNVVtg
V0t6xXDH8I8bnD/bODtBYkh9UNSO2TtouwhUu5ENkq12tle2jW7niq02DGDuDghL4kEVPHVbCrRX
O0wfnUQhhBtjBa4+1r+aU2ca42ssEwMWDgkKazjXLJyWz+D9b0zqr19WORMGyvtI17VWPjNtNHEK
LmWhSpB2l7n9l5w2jvfd688q4Fean6eWQuX9WUraWrTtpte4LQd4s0WEhxJ50AKqesgDRB7c2Gu5
wv6f3aU774KkCLGfqKkfLV4uJya/r33G8NEgXjqoDxv99fJxuiy/0t6eaIsMYb1q5OEzYMfVVwa8
tdfUUuMGOiT4tEm7cY2djunPO78HNJaKokLdV383FH+anRs4wZaL563ywR1S7DjTQGuJsEdtACNq
EfZvU9F1ZMtFpM1qRPqCLA7D5GQigEc/AvqUESEVrNL8/4O2H1+GAhbcVsy2438EVpOAC4y2ahka
xn+3HQ/o+ncXCk2v99ufBeVXfqsRPTeo08LLwbfL/AfzygRLHCKy0AaNF5sTtuDYzeZOD7fjqa3l
B0j5bKSVcJLjUjTzb7iYx/figBm1yExQD7Pib2f33OMjEX8MsO0XSj7HZFJWgJ1aJ214ZWfOrGs0
kwtOxEClR9MzrmRUANxORrVW3s9sBaRk0mclw/1PNCeVY+i7TpVUCa/HdIY2qTynRkMKP1DdTcNt
bw1BvM8gfJkbmIt459vahBWsIbSJuwbNAMB8mrZuMzg1rKCqC7yC839he/sU7GN6ux2lJ5dTDKKe
E1Fq6a34cm2MWEAIz7ae0hAr/QVac0FOPQM1dfnkAse5umj3M46xK+L4w7vmV0e/QVENqTAhWJsR
euwvqMiqb1E2URY473WOWB6H+paxW2nF8+p0Btzz3DSJ1hF1Y3bCtREnxjXGKRySJqQe62jq2xbs
ViZ8RBhVVJYlVv/efscPY2eTDXlLrXc4XAJaPACYhPH2uWtrWnCpDYrcXOUFrUSlDOvZMO5e5cHD
0Pah+ZaXkf5dSk74ltlKOVnzzss3YjHIyZVJ77KinHlrIqk5uu8s0LyDwapu3+2zVnB3K2Ti9m51
tqAFub/9asw8kb3TpDC11i/B1asA+cFWYPFrxEtjkyPbnpUkGm+zFYH6Xo6+bhV8nRpuD6foPFYc
tsa8HqEs9NViJGzmo5jlc7LUqFcHmg/xDYLu2C9qVMmyR0fOEVzPWqpgTlwxQoOrbz5ES/U0S4dG
jkg9Hfywn7YQMMGlWhWk4YEdsRKQFys1oux7bzqd79aU/y434iytlG8dILeYMNtfvFr7rUzKV1DE
OpSxIteMkGADe4HpFr19npuvim3qZkc+qO7mn6zLSd7Q86yZrcO5tbEOhh1cv3yYOZ4oIwA7AQlY
jhFcFongZlKa1cdj+o0blfxChrsUntmpmfckialxown0dszsSMXsY48yQ9hbNuRTB2E6COWoNhJn
aDCFRw+eknTis3DrEjpBkutKo7SIoml+wbmc4+VKm8fThdMjKLnTtipHp25mrWG5nh0bK13BnDoQ
n0nw37itgUElp+zTcIFUn0EkUzHOXU9aarAU35fu2lWclUA+p6sTkwUns/ePHBONHHpYMTkK7Dvz
f2ja5NKmbmmEAh0ijj8xhC9y4MBHtdpv8vf6wxOYXmYYBQtHOIAXDClAUSoKipxdWLewmq+nEbl7
4dYgx6nTm7gzLgCv2qysxRRfyjsY2RHQDa6+pA23NkKsXsPaags1j8ybB8nftnJHhfzQEolXIrGS
KGeq8lRmCe7U3dX9tPyP1ufEYZbK0R2A6n2MRbryU5UshR1RK//P6brAMuM+cbLsWMONFFudpoqq
fL8CAMArDrD+PjA/QIduzgIVK4xf3Fv85RWfMg/OlytYG3c9Lqey4GOC2mlW/Gg1wsdP830Te2JW
NB6Ml12U/adb10Yy2IbFhXzFEc0rW8bP2zA7sPm1l6umhkjTAgr9636XoXdCaIxLWl8Syhvb3A+T
CE8tm2HnnuOCoXVKw12ttgzkPKpXjfayJmLOucyHpTwOqlf1Kjti4GZq9c5CdUwjQ6CctFzrplEl
bnupul4DXXlE5jN0SdckgDojpD5xZ30C5sohuJ0wnMZpcebNQC9WIlC6Cotk0DyiBNeQppBA0jNR
dyuiKjG34STxdsLTkzMmISD2jkPLI1/ak5AhXt24cB6YNf9i5N92Z2rK2icW0/wGle6AM2kryGBv
zhq6SFrbyQQAfiDEx9HJ0evphe0ro5sebooujWNgeCpQF17CFfslxho96eJRj3DyPDNkwdS0bdEa
6wAPLcNYvrL5oH5QkAwl1BylSWPh+boUZt3ukgxtCsAz/nGP00T/iH48NCszopsrwHfjS/2LZEfP
MShzlJPIHFO6Op1BT/bbGyLKlozqGddj625bKhxuoV+rKmI2TVkiQz9xwbN9ZP6t7g1NFgY9IQa9
GWEH3L9w6/PPJesdRqCnUOWtYi+z3+bREt+cKxTei2iod4WdNGbGUmekzuvhZjr7+uNwtcWNKnmo
U9pqxEhxI9o6+zVSMDzUFjZ+3eCm6iytO12oo2Cet95M5agRodF8AgFimP5F7xj6tdFXOf/UAYol
RzUm68WWSOpYYV4bVtvloM+ccZtrlRco16WrY0G+h/XzX95xB+goQ65vh+cEVZUSdjjWwDlT8kLl
/sHbYqPuX+gEs1PB3HZIwQI6/HyT+xWwVy7hQIADyzNrgJLtynXGUTTajAHElbrl1Ci4lq2526Gi
L7xvcO4N7DuK9p370V5JBgVgywtL7zSFA0c8pMLiHNPD9fl3vW+9Plf0FzLMX1qhtdqCXl94nHL7
8UUKMADiON/WcCnMF2oApgPZInGcREalt7FKMd0k9sjdJBqvWxlAgc3iYBmhyUAPvdO6V0/nV+nl
XUX55o+8YSHX5DgUqQEhebYb6NKksl4RYAIICjtCczE6JPwYnUuQQldLBiuDSFLIAS2L+jqXtZZQ
wTvif5t6vgwS9rPf/Prr3xA+ONxBu70bNTOMFrXop/6J9g2PNsRglR1PBS/HdN7Y4TOpOn3rDp02
sOPTDPSA1WmMzE7ZEfZBTgFLp1HrzxCa2tE0to3TC75gqUz0avNeadK3otSXEDBFirMQIejXmrBk
yhC6KnLiXYvqG72vw+Fj5Rq/ypQDYOUmoN49zsJsVYh+oWMwLCGZPpk1kq2ccIxovTh/kshglHrL
+HrtRtQILvmdJl05+gwYPk25T5yHhVTuAa+x41pWDgG/fMH73gtNnKRtAKLqNjEmbn1xwaFgobxQ
bLUP6PfemkopsmVWi7rUHHIba1ujHK/DEZXOqwfVKVil3/l/4ozHOUV6JGgwbgAWqoOfbkX1uRLi
Qs4n9U0ldOWMDYBAZKD8RGz3/HOwkAwx3appqgqhXxwWpqJrlfMekMH8uGH7AfbBrbm6dCjNZeYj
bjsnZ8Sgr+jjBdsB2Vthz3EWYw1E4Kbi+YHdhEtr/9KmNrnFmKqdBsxx/0xjt+Uh4s3vdWQjVc5Z
Vw8as9k8SAMoce7vRYh5vcW3uBgZpGzxJVAzKRjUWLRP9t+zqWBjJ5jk/a0lSWGR0PGuSz0vjqID
y/crrM0zQxn2GPuSF3RKX8JHRLW1YOzhssv0irY2sQAx9OVOCmRUcXjhyVezSsysEjRV2RR7UEXH
YfnqWflTtmr+wLDkIwjJf9C7EuQgGWlz8Ivz8LKi1lpVo3xGfnpQ9q8+Q1AW39Obf3ZNHbDN1yxD
Sz5ONoiMzmok/slhSRl7F9j25HD6k3uDbgMeqBEiZuhluZDQ0+apTL2Ta+jZhpipoMHjuQxhSP6B
m0SrndqfF1x0J+gpk1mykTzumAhIQYLtFFhJ2NuOoqCBeN58WbgW0c4vJVsCg5kzsxlEa0ru4BpX
eYHmb0kU/rNf5yvA9wWQmo4D4gI0a2gmt/APeoR+ifKbV3aAgxyrX7F1vE0eY5bgiTwO1ApDu9Nu
A034HGEz5fuX2EIKiockDg5ET5IGxclrikiOMR6Ck3K27+VDtoAI25ShU49rElIUNAnXzzIkyeqr
2VS1LAFumJo0aCykKx2PdiFQh49IQXMHWvQcoh1wHAt0ZbXrD3Ga68P1C7eLJ/I9cOjkPpmCBrvk
SJUw3HX26qIfqsR17Lc1/GHHeAcE7FsvLDVgkjn5ANw0E052E55clniJPiO78aFT55+Z3Xn6tkZ+
U4mJCZCHPexQhzbYrBcuUAbUZi4W1jFXFU4kgkofvAxqYdXdOuhTwMMLkS99MLr4dB/a/p+ipt4w
7LIAm1STkGZUSDfY4lMH/iS3rAYK+sQczHHVqXqCwmeIlJdpl8kH11kEQmGxsZNbGNohP+v/3w9y
H1nlWj9T34lM/+ZU7c23MRv50ny7UgDHjLo6+sykzfW9OkVgMvIRKfERoE2hIKPbLQATtY0XfiF7
q0RQTOH5OwddduOecVzvd/CWVIRPrlqXNrQs5Ac1F1nEHSFAEnR4geMwzMr1RoetrQOR9Saq8hSF
kX77y+UBJlerIK1kx83s7JMkVva743q+71Q74FDDXJxhqy5YOTP8SW5yKBfbncwYAl37wnNBU2Nq
DywPgtVaAF0dNP74ejeMDAuJlp8B7fRdrOcF2OJrFhqdZQj7LzroFnFtwH0Xs/Nx66CpjAn+yPzD
juGGpsIZB933+szmJJSqEe5OmRNWe0MbIwe108VZR4irRv9Gij6kdhvqJwODYkYVVlslnmdOwLJP
IxOd2mBol0hZMuJJr3FhjgXYnCcCgsjGuthg4/4IsGAs5XtV+0VgbDx9+oXW+yelZCIs14GzdJXA
oVLQRHCzOydOW0IPceoDMhEDrnv+xYHkpiWYVMJpdAAzJ9DzURhRGEluCnXINS0/T4yYIgcZoau5
1jQArHyylxk/LcCf2iQeAW0PFA/aifxeOSkMMqmeiKWaWsNow+rkh8oZlX6bsyzcSxcuwxUG88Yl
8SwfhSbOV5wQ12cePRpNMDZSLX3xKlrgzaiDHwwpQhPvFf4swNIx8odzSN2IGFUjxfKZNLRR8yVo
FoYgxR4Wtl98m2bmE4L7HA8L/YceTWro7GzaJey1Ht1n5/1IET+gyiDS+horfFrouMskeAwOMgZu
GMfvAW9GpLZQcawc7GPjgHNxtX/dDdRx/YrvoYHegb9p4lMDzHs+F7ud9Yb/AjHvRHKmz4xn9OrN
1xDcVqMiFY7xrrbws/zqK7gjN7NWRJzx2Im+BR3OAQxxd3pxCkNU8r0I7S/uMKJlis8I3N5u87xy
td7gtErIkmeu1+gVN7xtpljuEqGZSZxK4MMLaMbYyFyHTWeDK2HWNZMMQdpXE2Y2CBOFF3Zq6ec1
MYUYLrFhkdrWqvZg6pK7hLaDwoWjy2gOs/VzPbqcF8MGUhwjcZC2eyTtCaOYPJrWeHok+XyMKtC8
dQHX/LEwnYcjt6KvAWPjh1AVTL32CvLb64xWYXiuQ3+mkJQiZGqv2XYFNTr2ArAwB0e8BJiLEdzC
0zwvFh9TDXovR7hymUHKvgZuwVITzi5WnHEqaetmUzqlJ/xMVakOJTHI/pW82f8GQrPipzNO2isH
XTRmnzHzRGaakc5Igt93ZLVVkSTjGRFd1tTZgnoQSrRE3u90zk2IMsAazyzgbmc7SiZHUN1hD+7n
dZBGlnRE66mtci/g2V0Fjt3p1M4G5N/Ge3EghopnzmCPErHdcbJTs9oAvH68q82x+G04JDpzQfTb
C+y17aaTUuqiRC6sdi/Ld94L7HDrYGSkZLbPes4PpA6Dn5jAIHOvdcne7zCirUSB+f6l2Utuo9zR
drUTQqqVi/goQ7Jt9hOLEVj3m5vEI+A1QPaaFUSU+XSegsSviArJ+dRMsUrXn4srKXs2WWWOwPQb
WCP/FF0vA+UquDuQ/DKOcWVhQ8Om47ETzS47SLMD3m5FjHBpsaspDC/TCzCH8cIDDMWAJm7FpUxA
KWP8mesjK1e2q5zdSqBECNd3aVFK8JK9QLwcvctNrN4qIUXDwJiiwII/bDawaFYeZNGbs1/jU1IN
ZtltTU6wFU/5z3IQtheHpP9EokGDYgMvsI+/LzoW9uOk1TRlvdH19Ey0kG9CJG3JbNaQXdWLLtFC
/uMuU9UqXSFvbwFxTj7mE8mgFMuUuXwhbkS4VvZGunUZ4DqH8DNdQ2v2AZQzlUlBx++cXfOXfWh0
dSVbmkAxPVfnnKNajtWbjO36vJTekTkDeyNuOJdrzEgTMldqthZoToX25MPwV4k6dwHgSCm2xRjd
5CrzpgByl4ODGhJ80xeTZaW1cCwPVJvm6g7k4wYo9jrlm7AQ8a1zs8HaUqNcs//99fzgg7YrcVkz
PRI2VYXjNegaEgNP1d4xDaUJNwaVf6Cfe/Fm32vNnIU2p8sAX9cCyp2qpTQdsVF47XMQMmn8eInn
RwU32jGItAYo1Nv0dsmMREKBy0P37tqRYqq6haM/gjYxZ4RcLTzncmUrQhxNgeX8MUC5f6cMOtfU
9q+Xg0VCBspJwxQZDBAGkx8hUri6k8uPQLafx6HW7cBYqNK8Eqgvqxi6qxaCX/xik47myj61KC/I
ZcwLbXIL9Nvw0VtmHA8zpsPB5a33/GrmD6O2H3St77uto9+YQE7EXEJYrBV99MB/h3xt2rwAOwFJ
0RlNTcU3ZPcV00iMJFkxx2TIs9sVmt38lJBhqtlkpRi7yorfNPwlbW0M6aq+mmlMgZNmdBc1zI/R
AZLv1nC7x/wBamX3DCu4S2bvDYBwaQk1i11ZyMpaz6W54LI/kOuZfKy/2WAh7BaoLqLkCH8d33LO
WtRxAxqI0QyaPgF4Koi7WxqihZ7mJTSK6FFrxBTKBVZlKuFUoeOYr99IRo/yw5vyRcIrTxjfKYOv
Q+GDGQfl0QfrYPHEugz/XbTqpylJ9WjvUoEVhm3CnOy2BXURpoWvjRHsdd2zsfEA6D2qTQo9jrKc
wX9FxZ9Dx0kOLfYqdMMNED8O7od9PB5Z+x+uDgY8xqNZYkx13tvw+BF4vluL+2GQVPPDqsPhyAO9
1UbUWFPLwzmAt5aRPZvWQ0m8Q9ybNkWEovNPqExag9UVP6h2ZxV5oMt2tqfFCLVIn5vEAtBzeIXy
KC8hnm0maNFBFCcIs4c+nHu9rP7qz0UM2n4p97S2/ZYxGQ/pqvNCVtt0U5gLKBC+eUp7T1x7rK4Y
Vc6ip0L0QI+s7xD7byzm/PUN8UuaH8HdwGmpiR9q0lJpic3QnzCFMk09yBN/nJxgOBieDjuzYUc7
h3hZIZZQ6nIWfxkEIvzVBR3BiXUQ9ULTRxN/wtR+vJWuXPlgXcl8AjT3/AqZ0Fj1n2ydNvYqFOR4
EOqXb4j0GEMnnRV16DrsTajCm6teI68J8fsl/e5wWb6ubWYci4QYMdp0TrRAmTXBsbONQ2XjyfzA
EzbbHZ8WjGSrp4FANX1JJorRv6m/FG8SSgWhTO+x17I/9iK1KFDru27UCm9inI64mWDl+Pw1fkQh
0zk8k55K2bTtdll68NjjGHnbxCbDK0jPT7Dep9TbSJacd6Q3foEDB/WjMAKp3h0wVlkdWltBE8f+
YRqwJHM8Mod6CTzMvwpvmLciFN9SA0PJC+Mun2hRQv5Y6H+N06dcUyzaOxT+rM54Z9IXiv9WokEH
ybvgZ8YoW/98KX4e6/d64lgLUM24KXI1vV6qbM3cKb3ivLDOAKztuDpR4ws1sYf0NBOzPdr9FfVI
PypvvCE6jCPv9lv4jgARFsFhfc79atpMxOXpTkCdjVumbF36ownOvSDu7FKyoLyZakn+Qgjy41MJ
XzwUC0RDk8gcM/EsPOF9HZteLHjQi548Rfk1ImpUtxnJOxZHY8VtZJfeu7d3Wymib8iUuuzzeQOO
aLQDsPsjkquZphDXLViru42BzESEx9gaf85tFGNzgxJrhHIuTypoyZMps4lFeQzbsyPMEMI+R12y
wCtjjWCjAjW1+fs6iPUNNd8vktQMFgXWX1Trt68cpZBZndPbN3WrwqR8QGBVlrhZ8eGu/cnAUr9s
hgE/ZhiO4QuHxuPXIfXrPgLMTapz3010k/AFX46aACkssG0FXZTeHKDIQNVJVQ6Di1FRZhev2WzR
ZoLydndZDgxUWppq9XC6Xs2IUbRyIWLGF8mKtGLgLv7YBFmS9eLf6aqsIIcNUgmDUyYuJi6Qv8ZV
uaIoXKF16Upj3X9jGnTBr6XKCRhmFORJMIZfBcwwlcJ84sN1yvsIoXNQmxoutWmcubY4T9ycIlz+
BaVfRZQJecj7zZDh746k8zdHd2UelPOPVGVlMzwVZnoQCrd+wApZbFdNng4cRhcYbh3LPkv3sMX8
iMXjaWssXU9EhG+PJFD/u48m3aWRGoTXw9HG/wwAcZyj3pAhYbL0Gj8BGHfo+St8NyJmhTwv/7+L
sMIPY58LwhwDlGy2gTODkVFBGyYaVBNKpE/X7A74h9WbyRr0qSCNJQWwdz3+OO99mZZqRRqWjOAZ
ZyETDA9iIZ+EMe7JX4XlOVCP1eGCtyCXSISRBeHwNSOSu7qsxnn5uZtg3IZkqlag3CZdNXi+SYiX
DA0u/n5aHKtDmSPnXGEPSBEeoELikV58is6ksUCmoTxdeu3mB8QytHOIU05bYvATKXQMloTwTzR7
a/+QhPezI/x9SLzQgw/Gl3F+bHkY/V6g37hjXoJEUoRg1lGgtWNXs7tpzu2/TLYPgRxfOzwpuCfc
iD6ua7ycm0qZYzsDBR4z0eTFXNGOhp/oH1wPuEaPYZXQeSG0vf0ShzRWvJ/5EbZTuufqI1YvkyKQ
IF3m53T/O89ZzKPLbIzK3BztUiUNJZfp90aJTzWv3KZH6lThBThuoqU6ftsAZTe2cgV99E+fjmdD
WWOIYW3VtI8dHx14D9edLPiz1QnWKwQxJXGxsx8JafG7eZtTsGEDk9OPx5JmpVMOU0vX5g8/APtw
zm+A189WPt1YAuwPm6buiUhLsM/vrFrQRC1GMeGBosMayUYgaPN4Awe6hGkdskcLCwXpiZAEHk29
EphFAzQJP7aJ4vcbCqXSFpmWdu0CvUByIESdaqD/RRObSs2jrWxXms+Q6I3UhuKYuCHlLASoiORt
xkAnQejj/BK9Y8ckA6jB2L4NaU6mfRegT8+3pfPhWAfzjTgnmhE2+P6nwo4UWiOzHwIRCGPqryp+
HJeFpW2NyE9dHcw9wbBMdV6GC4VqYKuYEht1MxOE3cyg1suvq94+rktZfwE9r8uXBQO8XU+sCvOv
dm4QVzyWUXqBbY4sVGlBP/R/hnysuuDq9mhJ15L9FqArfD5aAqg0qgF+RjEtOZyhuzgIlnBvYUSv
mdxJ7shzEsYKRTr4zHJ3gpCEppSZkve7YwRwXm1CKp0xwQW7BFPxE51UWrUOLk/oI+h52170eKQo
Rf3lT//Dy8JvPosjb3xQy9w0T6f4+j+32WmyCi6PE30ESphkEG3z/0CyXsMsrvnuZcgN6fuKg/CT
UJLt6+9ddk1MIZ2brGZp+txsMtEICaYEVBRwkfCJBAsizpnVm3mNCqRgyz8PL0qrGfvLmw3ww/Ux
V3OHkoozb50jSaQd8DFxte8cQQpGbANAp/frX9Gh83M4GaIdny02fyCYq3oUgIafvQaOXRLgqIC/
1Z+qv8rgq3CiKzBwnY6Y3+2pWaA83Hl0H721Oey6q51WhDhmoIV3qP9w92H7rO6sm/NQwsolqEav
TV3uq1haDGVwRCrhsRLatr4rYrfiGAFcDzzfJHHWi3oAJausHXX7hJ8K9qeCdHTg0hyL3SqWrjXB
YVoZklqZfT52/fVwdaboVkRJybTmcOK18FljqDbvBtSvEcKdwkOAjWstFDDWL2JyHjIi5zm2FEl3
xIeJ/j+DpUyVhYc6Rq3WHZt7jUKfqTaBcGRExOTup2JTOPS/ZujwMWeBhhk1MScC22//Vqm/ZMVL
ji7bdfmI5qmTJXOwGOlAr0aZq7GQV+HHWrYq1diq3bAGfwT1BQsiW4FIk1twoKKOosImZ3kB46n4
1cz6GywSls0t8aOJXMo+1VC0aZH186ULrbWUwVSp554dy1Rf706MCQoSHN++oznYXJ4Tx1oucYDl
OicJ17KbBYovJps1agk1rZM/Ud9cgvbJQOpzMRk15ki3MQX+exfnfslDrmIC4T1ZMeYzGzstsxK2
9dOmWxA/N7kiovjapitWL3ywusHLWMWn9Uj/Yfm9H4m2W0bcZEWT39g5NZctLgnXKD/Y3EMKKpsd
w51mMyyZV22skWVxJxZ0OgkT/YlTvya4sqPxogCJs68NkWaFywIqeVePNHtRoXYlF/ACDFCwYBqL
2hF2cLuMJxqKbEahqZERUxjZJ7dqTo83BycFjEenat/qOrPBrM71B5GIl2mJoOEUWZqSjW6k/m0W
O5lG4riSaSsgmv3nmi7ADiPU0OJR6JhwIS9Er5Vc1aQL1u8MvnZq5RTNPwpcZbkG1CTmmVy3eHxA
FIjQP9/u6r/wms5Li2RnCjFL9+24gksYflWidOvUSK0RqUvnyQJ+a/Db8KqWNHQh6psz6wcECgxo
qftWqoXQmEM17YS79WrhnEOlZwkhCY0gukztHucqlDQ/CGN742kV9ZDPnNH/eo+BDCiSEs9WyWP5
Xw0jbjj1e5Al6Z5zsp554Gvq8owz/UbLleTPSeuOy7FQ/XxmXCHHRNjniAANyNo052ZwNlVGDohC
Rv3f0iB660IoDbKDOwlxO9bHRu+SlmDtIkOCB7x1V2RSHEvtWe2CydTaT6/C85UVbWnuT0Dj+wKB
XtrlAdh/ifnqRgSasIYneZTsGPObhHVwPyh6uIy5gkOQmocy2Nq3SCutl6VlHLbN2AZDbL4Nid/v
T0ttO0RBWFTzT4QoFaxj4BUcVxGH0secVc/KyElPyRv1nC9mHdmiOkPrFNZEhbURN6TAg43zFqxu
FobKDZ1iK/n8k6YOpt4zH3rSwEM32bzFVecgHcg0m8JAGTHgX5EjeVefeKb39Y5V/kJdLAQGoOqm
mH3KHm8amwi9ZHBN4CkNJdJRwtE0F+GyRViEczO67IX/mbzB5k0m7jv21gepDi04zFISANgBZqB8
jxJE6Otd6rAtV3NUQdhTE5Hrw2l9XWnYADqYHEWsWElgNBwB1AmaSgnoR+qwXxdfJWm35uL6gYNT
r/czvVNMHRttqg+NQSZ51bQkF8/lIGVMcqpQg8bpr12q0SPVomi+eHKNmuPiDDtyetZsdvBNvPrM
4eFeZrSfMvsOp/YwEyXFv6+0f2NTJjefu84uq63vt3dB8QS4gAAsJqZEVS0avcW5rmgj8OpuKoW7
sIy2dB1gVZ/kcKMjBUkyV4jxuAGjQ0b8foXOzekIv+m7C0mJKWYp0wpt2G45vrCDcDW77u/XoNyg
oJDDJwMV+BL1/513p2DYrz1lEj/5X7hdcBp9bUot4Qv6e6jnmfbTjTWWC9rd31kFxEgbpz6nWjzs
5Fq6WLWQJiYd2TfhQQ3yfqQmNmOrCFr8jkakn2DuaW3wGhizrb3wOQahyFpWZPr7Pu6c9bg5NiZP
rnwqu5eK/2o4i53CnTfnr2EBTooIjMoArWME9ISLADO3qL/pNFYcTQgEWQ3w0uLpzplOg/QjjoFW
W0ALcBu05i3X7de8hFK+yVhuQGipw0/5guABPpLUYQjEtqLJxMR18CQHLPqvejLrjqYJCP0rDa7K
JQU/Q/9sWGeddW8V4DawPVMDtJa2WPD85A1SMUzUpcaMq50Hf3GTwvpieC80fg9VQn6D+YMFg2EO
mBJAs6FVJ+S6nMudw3Gh+rLmPrPgROKg8k7aL269b92q7RVLcAFs4g51mGN1k86IWN7enPDS3Lyr
LljbNRxA18F/TM/pdMqcNBIVOKyheiT/PZ9AvxrcjcYKsXF0nzsMG1/qfKwYgfLd+1P13OzXx9Aw
RlDCHd8vpWbwh7lRMfPssC0CJdUATmWcJYlcdc8jTqBaeyqzxi1tKdGsaVt0ucYkKLmu70a5agwF
wW2hGzPdAtZnS1DB9nwjVtB47Sa+nNPDj1i60yhVse629eWmLGKY+3+rKagJ6hrtERE9qzyo0EpG
gXbFv00ufLG2jHOYYzLyGFpvcLwb17NQ6NgLGRTCFQfgb30zeLyrWBfPA1HONuG1K9qDZVrFLCTU
vdWVfpZk1+mmcFgXLivoQB3W8zyKUDDsgYJZQS5cYReBzg+hFnXSWMnuE6yzBfL1iXlfkla5l4Rb
XQHTF6lig1wbh2ISh0MNbxxILyaXNGdGmo968Wprh7++kG8jdHPfCoMlFSfgKWnmGmTkIuvXuD2C
bqKOPLS38cpG/rF5uKKJOrqxHbZ09MG5uea/tplROGYUNdZRbx4Xq6TGfuoQJYwq/AjEcuc9Xrcz
cqngzQ+MbJpiZKIRmqBVlv/4PY7ed4KGwLeSAvAREZekp89v86pHa1gVF7klKIRh2T+1qXyO91Cb
Vy044+DlnoVKrMsrWJG38DOHa4X7mXWsq0OMHiMN2lEOWoA8ZSwrI3JhjOpjL/9XUVu9r6KDCmE1
4apLUHnBuGRnB0bggkXMaAKdfzGlw3erj0QO73LxFtH4pChmlDF+NY6KNl6SFTti58OOBnKNk6yv
cP/VR+IUMjYnMgQDJcE59KOyLNZx8S0zj+5P9eUJ96VCJk+XEk6LWAVC/YD7+bVXdb8Ik98XX/oy
nZXisfxQ/ZH8N1Xez2VGk/sWtzQ+23cSLn7voMTeLHlvQtIEQ5Wc2qiyJCy4Atr18p9NJIxjogOu
peh7tfeCjnTV04CRwJLwYCjazUHKDxd9F6PUpXL+qc8Top/u78voDXrCXsZ0OiYpRfkJgCq+RgTe
1b8pU+eRN1pnTCnXaBzvJvxV4aboJoeksvpDMv8lG5xqghhDPyu9myx5TbVE08l/dmSEzWPxv2BL
bxIZMFwxaHnYWIgEQb8+xiHR+7uS3nhu7ty2t7bqvHOOVPdFA71aNKegI6Tl4NAf7Yc8aV9Unw2M
bNWvkqZUg5ZXEvR9ANgTicsK06YUVdKI0LKEps79vCs54yQYEx/JqRL1UVk77b/8JQid1bWv9jtM
b0PuqVPLDL8vtm2nZWr/8B3wS+sgjXjisUvZG18hxVKgat+/zv1G6iII0a8AIYPuEfbW1UyxhhfD
AcE2KtgQGFBRggdIrCQRMj6Xv2D6JikPd+oYUiBQhgiPIjMyJxKJK9S1NnVBRNX/dGS3G9rpkB/v
Fbc6NqhlNVbgXRHNFDUZA+96i0ubEmAF8XZBN55oGzzAc61ww7SQuz3uyVITSyMQ/DUXhEJ6XJf2
CAB4MVlkamsDjYfkGYKpLI0gp0g8BKtaDfvg9MxM4SvaPof0dxp3V5IAGL2okMTfWPCSJ8Dq/oKA
Yo+21myGIOj1e/Vq+w9WzxMPDbwTBEoiA51tufPR57dm5kdNSoMYAEi8hN6VkixffgwvTOrFFNR6
9NUS1Ph9QSXsdhsvIb9jOjaKqq3cS2DR98E+ibxhZ8834SZ+awi1Ei2JkSULM/GG2j+emeMyDAMt
wgotLOuIgnpHNftN9WIHRE5YDOFAIcEfxzpnnjKj2QkM7XV/0Nrz2xRnLyHkzYKmbmq5D8RPtbUz
X1J36IjIQDf6lHnF4H0+P2MHjxY0tw79fAEn23qXiGlft7uObTIk3i6GdDFpNJTqVDDaR+RdXELm
0zvdAWn+9qzmDcvDN6wiBlYrYBZ2BwxIcY30ljDBfMi0Gq4UokSU+QXwM53PiB6cQZGfMNvi0BpL
oEv5wBP/f5EvHD5181IUzsiuSQI6kTtje12o7pD7STV/+XTs5DN8IzOhZwtmUjdoMSm9ydG4rjrH
+zuWkAN0BbWapUcbKjY4jQvjC3GgPrEMvofEgUjCs+GFSD+dD5WOSixMPcZWN2dnvqz5qJh6MjxU
wewJ3eIP1BQLBoD39bVUGjQ7uZZRfIJeCrU6OmSmzxjeUmOfa6fE/Niy9kgPgSokRk3EQi6/Elwg
ym+TVg4L7kMnEoKYR3TSybyBNntOMfIsrPwCFrx5cQ4SWBdEcfkY4176Cg6R9RHe7NyXA0HFxw1e
kXdAWGZ0LawuqvYWw3SvfONWqpcf1X8ZbYgJPZ4qA2NDmlhjthijh8q9CZ9FhFtnPtf03o78i+q6
5TOa9WT0nwB5imMG378dz+/BlBlXf3hTygdDiQnx69nCikb8OvNLXAxagS6g/L0c428J45OCXSkU
S3ZaJivUm13ziJX5PDJAfMA1/mePktwKovoLQ/5r6AGJkjO+8zAfejQc1PjMABzCmq1PDoppvSYG
OQ4mHG5zVlTqzBOcMvmS2E45hTLnd3Lc0tEyrLHND4JAaDnUxyFI8yfVg0iBKly5iGDHB/ky2Ye4
cjf43t+0HMcXo8YpWnJjJ0Zz+QB0AAja6U+9XaNTKOSVI0R/ZQjCsg2aMfdf0Mpiv5S/2X5SmXr+
CgGSU5teVzX5gC0KdSnusT7WFk5ssKf4gIVFKtsMxKiiAnPk0FNZhG5T+uobM7IS+3WA+fkFpwof
6mgdpav/RDO3Ak8G8ND0A/Z5wmqTKqvwKWW6KJlMrmPIk7tCtKSbMpuG4WlSMuFYB3DPiOqponTe
eUcn++3w7arjfM6O/9J7RPZI6mPU+CTQo2gTXGaT6Y1MvX+cCcpcr1UpH1p2nyVOCOkDniQCgTcw
mO9wUgiA7j7iDCkI3rCSQCV5Oqos9toXmFGJqYgadWQQQtyXIKrEKL8By0n8JDM2df+kYulBfU/Y
TpuXhVZMm8RVlLNbmqkm4RsjrEF8Vl3DDJEhr4Q13qTPPPUSturQb8iHgKfGqIcDVMImnToio+qM
SzlkYq1ZqNjXRzbt/ptMAHIPdLMEEMvgSclvkJegM+Qvi7NjphFu9rblxWZGNg+DgkE+ohi5lrAH
2ug6kiR68iHj+L+ovKQNCzRHT8YNZBBGYuFbVqTVTCaWR2r9T2zHkpRfDefNLpacmWVCd2QEAc4c
FkXQOljDAs8XptIPpo9O4viyoKcPwsH1p4M0M2sv6cfJAoyOSsqse6NmFOs49a4p7OO9KPShvV+l
7y7W4LcTAetzOsX6TbNIQJrX1/ZKp7IV3iGiB4IdulLyWiB5nDFd/FfJzYmwSywlDx2/W4MyQn1s
XcvMniZny7EKkoQ9BF7Bk2+ebuUm/0ETtDRXRfHf846MP80wl0zXZ2pOpEEnJWhcMja8gIWOwxCm
rEmLu8tEzv5YzaCJ7Kqn3ZlyyWHXWQNfsSlj6ZP3D6lvSXZhW3Ux8PzFXb17PwgkXCajujPQnXP/
2YvZfh9pKd/R3FEdKEgduVAiYX/Qwdd+wAPTD48wtCmUn28tvRgS9YmpsDWLmKUhfj5sMrXvz71S
+fV8Gd8Mguu1BLOg75dHf+7cjQ/3dyhZNam10CELMpRSu21OoEVqrp5jd3z7iCDEGI6Q/b1c280b
VgasS6J+xtulZE+vUb/U3+X9mPmvSIKGQJbcYPdLUSRjwPRDCHIKNd2eAqbZIy01mdaBiuIgbMtV
OBtfuFEshdWjmDoo9gS6sR2lnLRvyVoY0eYP2zC1rhhmrh9ckfaa37GZB3WBonp02qk9dXGXAL4z
N+yz3xl02ANyqExc9lIgTAs5LsTOgdchDPRsS0uRE+J4vKqohsF0dddSC1Ol7AfAC6U5WTVB6xoR
u8wg0GCazbnX9VBAdKIFHQKHyMSYpgkEXK9s8WIJYfowLKR16NJc8u7Cn1pwiMN38SOr30lUIiNM
Awo4DJQ45mEnt8XqmOVeocYNo9dPeT+bIpEHfiGww9F0hhYJ2NVcYF4RmvjhChean9wG2apTn/8H
xY8ImXNVTtoMseFwNmQAupu+MC3MCf9w9KxkBiQtHPibCs8pY0X59TjsClyi0IPMrCZ8cRtmYdgt
CPG/9qmsPzcWcckFpFiiCHrQFI8FWstQKbxv/b0LMy2MGYQsJMyVd/ZxxhGiOlcnN32aV7iVkdBG
Og85uFf08j+DgUmpwuAOnxItV1XIS1fsHeOElaqlP4TbAkQpq4npSs6aBoFmEAQsazDq8WCDSA6H
dSv5/5C9NqFw5SN0k5XIWVVRewFGzqd45c7tDSf1SjfNJNjFW9B1rVNQtSyUanomaNIuqHOcSQE3
njJeZEHFj4h/Cd1jV2LiO9iWEE2Drehvos5GObRbR8OV0AgztwfbuNgA7bsweQtkdlBaYeLgzLMW
rH4qap3P7eDOHACqUOk2ud7aw9Fv/MkOZ6Qx8zVRmY2/FeWGP22U+uOjpDyNwv+yTp0kFzEyaN/y
R26FMUBs/djcWqTAk2x4AL1RcsZCaGo4/EP2yDswco2et5eU2cMOWcnejaactU6vSIBiWQv912ay
86FCGGVM55QA/AOQ8dXCGMhpDUaE40t1xW50/FEdz/fxxusmS4Ug/MY6vK4ka17jmDRB1K0vzvke
v18+2yb1/0Toodi5tmgW6qCSpqCHxCX6ZF8ejLTlOViOR9G8Amn89IlL/6fFWtawXTJVgARbxYSv
mQFgAY++rMjiI8WxAn5jvipYUF9X9LpLChZvcRnTOWB9t2+eYr9dqy4phJAijb+o3a4GF5MjIdFQ
0Rgdnf2/bB6w6VMgeEX5y4Drpt3qNBNsUCkO8lBYcBsomIHTc89kMJILTVGO+yRr7P9Acharhbt5
xmzo3JXgSYRUZHd3EleCeFpO4A4BjFJfRfTea3dqO+WImIJIMU+4SxbXUolAletTkmWkzGDyQAz/
jjGfhwMjeoPDdSgxe5ghXQ0I05V3w/r7wBZ2yrelTBpP4pODFpV+Pza66vKX3IwZXsJaIOU3K7Xp
kFavGnl9OMk8+IPZ+5UBBVdwuy4P/Af5iV83pUxd1HJ+TEdfB9WeV7AgN/XrR0GrOnrMtlXsAwHX
jlve7fcq4FSL2KZWtT1OZILAGFrlHefEZ423/6mhSO0rx4l/H4JGHskRrAf72nG6q4f6ojXXCzLP
wTn641SgYNYbIsmhO2JNNGB7tAgv7+lSK+JMVPusvYTZwZJM1a4RHoEg4bsEsO9RVhJYUxfypSXS
pnm/sQQw4u6njReymquwOaKQ4o5ytvaHwf8k9eiG+g10WUIoMQFqRkHotUiZzVGIVIK0OvbpP8zP
AX7AyLxpwWy7KH2W+nITkRCsTHiVM/UDos2nYFol+BO+16BCOBhMnmPVkWn5TvhOTsrT4jmdn5MA
UufJtH9yMIxytuxXeWxVHCewR4RlnSV/oiSsneP/UCH8O9h1OuE1OtslTtejkIoYpQ+lJCQZCUOq
0JYr6WiXCEl923K7kK4deSrypByBRQmGmw3KbM59Wii1kCVrTlgqMyYMLM020zt3I1GP1CqMAvmW
BAE48mojbg0Qzju9naPqjXG7SYAGZKXZI50+KOtwljbcws31gqznssIivxLFQBrnlA+xwHfQODB6
IgdjdeoRx2aYFmec38bu9I3DGZT750u++nWerbmTvN1xDh3hzA5wEArERB8iVIT5hccI7YbjWsJh
t/OXoos5CJbaVRaFnMOYSvZH4TSV2uMMlQB9FvkU3JCny6eEjMASyiw3QbPd4iBLocUWigVojq/p
wSfdWKlAaQUSN3X+OI+xx0KxJ8BiLqs7lQHwtA6ssceOx0va1a6skaNQTtOF11yBeG3HfIpvp7fJ
vexp7kUBR7gq7Yc7h1NB3xmEhKykhMkarj5njnTihrYNR82kSGwzkNenvZco5Bbg/y+Lf1JhXR40
pBwWaqbai23BGKtsIaQlaRlbK8lzBogcoUOXbYIQ3zgmwYGREClwr13pGgxUJe/Jhpiv0Q0/+fub
2qndwQOkpDPnqCE6DPaCDw20Iy5IOAGbC425pMDfxkvy1vMkwR/TzLTHJHrHPDb2Bq0Rd5TGrzum
7zhwgaKsqEh1WM4PhvQFg9SgiMAGcQkcEiTJ2L0obBjh/+a4R0bInEtnINKFTF3AWKn44m0XjNm8
BCX39k5qoTZMF82JhqxjdGfcai4LQSa2D6NHg9vzctgYyw9myHPIuT+pP2iCh5Z7twY6YMBXHTFz
i6VoMF10RqtldBO1sfwHy9r5MiCfUU+ibDYi/a0Dd4BXVm/PNPP7YTOnUHKfeEkozl9nKnQPUx75
AVAgLhQP1GoHLLLzGrSYDBftAb1rYl73I1I0Pn091SpK+20fvNuPSKkGDkssweH1Mh2yynTcrHO/
ZDhTw/9fFo/3sCn9k7rjADEc7jRPXTVWYIDG5e7/TPBs7miN/cuCkeAm2dubT7v64CxBYsLFBPWV
s/Ih18tpi7jGi+JuC8/i+qMqky1IBvI2BhlNPjHsMesPbnRGWIsM2qCrVLQIMDKInHhfcoYtlo/k
C/fT8zx6n2a/soDVWMdvXwQS9GLZidDaEu35u7oZkBrHvXHyhJgbtdsh7RvR6JmstBlP6x5e3Vj6
IRyxOvJnVVQBRm1SQo6JHlRZGxMnlNvXPSeynGPFJp+uVJAnHbpVAd163ISUMT6mKOo8E4GQ0G1e
yY1G2oewkl6XO3VE7mq+om3ZrFqs60Uk+hyKXbWYBtobBvX6YoKJvWrvs2whtJZgh/RIVmQf+CPV
50z6svgZZf5DJjTkj0BdgD3hHL93qZIip9T/jWs7zaoc2++EYDekkfrvIg0esrzwuHYAvfDN1vcL
NM6VycwKHElSaoB5sNDjJg5WwiWm+s5y67I+xfaeSEetnAoo84C/WVaQJUJTE6e5w4/D1RunWceM
FuOhVpNhqF2uhUEFHXvWI3mpUTC57b2UQmqpUyfyd/plWuDY3bEV1xZ+lTJOhHqXeA8JEU+pIyrO
PmCpt0Uh9U5CPLQrSfFBldTQ50/lFSipSJVK2AjEpRr6WZsDmwxxzs91rBru0glAUEBlzamA3cme
uSn51Y8ImEsTTUQ/NJ7xccL8Ds/Kq4BVGiJvMUplTzOzMIK+GxkmANnG+i8hA1aR5XzWH+cIC9cR
CaWtKBXb5AwPjlx3yasJ5oVxquDy3NT0THJ2ep2A+tGNCI2XRXM+x2Yn5/oYmwP89tG05ovgd5JR
lS7lVld9fTRLRYcJ2+ChoZqHUGdeWc6ridaxpPZ6hNbboPN7EMrQl8Q4ZHtFSA6Ss4WGd+m6HcYJ
Bd51DkqDdhZzvEsWbr8xP7CdZRiTJi2lONEpsbXax1L+BPTcBh3SCjt0Nfy59FvZo3YtFRFbab9z
10bCojB4iisBEWLrJGMbTIKdQ5cKRTLgr9nm1HksMpUt9ReKzAVCpCRjfz+/B4/kC6k+4DJGmUgm
18oCGs6SoGcIdVHh7y8smS/xnw+K25+YXwwwfaryhY2DDtlZCQNN8OKx3+KeHlzerrW9wquDjc8E
3B2rV1dLrHbDQq9gYJ5JFbNgwfyEkhOB9dssxRxuCF/i3wOTp4PL5zJ6kiN+9/w7NdR5uMdeE0Zo
+cfHQM2GHkw7EB3aujduysYErNd3eezkaewrOEXXcDpybGyRaTqVoElJNWCFLzKZXUPzjXC7UmzO
FQwADGYUBL68J52JDJSGSHugNluQ0fx94RoFtJZ+rPIQBZo3QBY1Hm30yRo4ux37YJc3g9e36BxN
9kH82miWtHk2YBUS9V8jNxMofgB0WS6V91z93n//ChepxaUfxTp9Bl8UG88vKieNBJy65QWOo32/
lH/+x4nLF1/ip6BQENJLJFKJGsQoc4RNVYnbpTatUQOsmz0FMPgEXADrazcPDrkZQ9TIq+0T+cNN
ZVhs8cUfS0vgZCu5q6w1iAmvdMpSM4aI0XNDuW7BOsbf0EOG0sjUvA3QtBh+dRsJwIiYpVqz3pGW
Dkfazgnh+V4xN2byZNq3GBAezS67d7qKuotqZmPw2kPq8BoUlHtl1mmwE2nic2t4zYjEKmquy1Q/
T9xbAxY7ggFvqepzZRvGNR8vNkQvUmknZgJTTOUJss6xTN0yosuzu8CKGZV5+eq6SMSkO3wPhwn7
arxf5v2J4MPTDDV/VjPDHKGXlWo0ZCTRm/JzTOTLuoCt26vg/DSG7tFBNurziGcLUxDlTJ9CrvsY
0T3nn9y6x+9SKwHzSs3oHS1+Q6zsaEXSws0SbHkUfJoI9aXdnv2VX6NGeIG86Aqxac9hFdrdcUV3
odvAuLHYcxCgEwf+Gu2AKYfExxxcZ20OL+LwJxm33b5e6VmXmIm+EwQsoHyEsQfJXUElBjveKi2o
vkrjWINAiKJlVzHNZBs8F/Op5XIGQAQ/cW/kpi+e0exm20lMdzxdpGR747H+/WY0/ulJaHWEWUa0
mnfzZZFEhroeDG4Ymz2mtc0b44AMhHWbdeMLQkrukBZFcq6CdRCnkZzrcL+n336Xq7KuC1egUpFB
hvcPQJSUm1h+IJY1RRYzwvg0FpkfpOYjulOCR3NsMsz1n6l6c9eRkSwrDh1OpihyEqkrYenHGvIZ
1e5Q84JF3ME/GmZvtHNhR6Cp4pN+RZEUIUk5E35heWOiXKCuNl7Bk5QL2uZRAJMAFi51VUCsd3/P
34YGxl2fjp5K3gZceKgqoA5+p3S1MUOvm9F2ijLItUOK2JUFIADNclCYi+kZUBZ5tI1L7T3Z/AXi
GF8uYq+ctXv/9KOekdLko02yVea7WqDtDucZvJu861YlsLue1KGRdUB0xiw3O2f0AUQU76fwHLfL
11dy26garOxGlZIdH883bwwV7CWWtoSfamETkQdEUB0rLTRdx6D7PG97BXOp1h3u+VLt30FHnswk
O1mpm4rNT87hIxAmeWvup1Vd6imviRyDMMLU9MSKOIJB2UaoJpw8BMpEYBfMuFful/Li+m8eL/ND
oyvJF68lpHNCJCbiCXWBnCmGAEHHDi5UFhS1HEbHF0VHWjTbY1ZuDON7n7hZmefW3+z68ZG3JpVP
whoEjUP1ELuK6wQT8JgYd1QP1Wn+jOLRQtE2m/Q5HzO8Euhkk9KC5JDBtNp9V5cA2wYMmtuwivkV
KtdLi0Y4Ll+foP9q1WGGR5dGk32JzI7OqwdKJi/h0fBmLNxkyNVrSY+YSr2HjwRB6BLgiLqN5Y8R
WBVz8BntTLQttqWfw2QoCalopcrrh5B3SQq1wVnP1iZRigalNOz8MZXvkmElv5cobPuDxlplOZV+
Ji0Ns2jJaV3NgBcdUPDWhJaGK6Y7U/KluwbU7UuJDiaEe0pDik27RELazaBW5+2ROSM4RLrxZVU4
iSmHkfzOk8/lJLWplZEcI5S77r1zxO4Spq1fL8RhCReSTAT+3UUOIrxPe2Hnk3ogSPUdCYxK55Mi
hh1Jk3aeAAjO4EiocJrYk/NhdTgLolxHnO1CB7uyean37NJm9sV5koD884Pez61X3VdZqrQFa/on
0wA80vd+WceXqwBn/AraPg7e6jYlYkUepmw+ql9PowvTKado2JZPkurCLZsfPwbjygMyn3ZCrSle
B4S9ZdWZLo9k4kaiZDzDfQf2YCN6Tn+a6nfjVSoxETbceZZlb85sSyYrA/ZFgFOyzCK2qH2D5X+o
4CHJ9bnB1td2YFHsELuD5GPpeHqGkPTF6nBhodnnaLKWZUzLOdamUoDUsZCN2eURG9zkCP7dfIUG
Idhxgto1lwqFKi6UkIKWenUY3l4fRxuSomH85BPCkRYwvhFggAOE57SdGD7ISfDgP/RMjxZtqquN
x+lkLhm40AGLRNyZxHiwCE/b4gD7t3PO/gM9e0CM9VlC7sveIJ+MXDgYXbqgSmpDlQBp1zf0hSq8
Qs/Bm3NYAQkjIO15egLzMg6Dw2x/PbQaJ1bNbTec24W/wHRweKMkXzUZhZ4Q1T+NeryMeB+uc8On
xi4i3sq9oSzHI9zd0bhBNQDwQWh8nS3tH5Nio6UhEx/kIdyRlGadEZzkdTiiWdwPWFuEHVrZC9oU
Mha+xfwc19KBgfD+vXorkqcyP0ZwtkrOQ5NA1ycMf6VaRPhrn4F562RYb6BMWsNJr6Q7TXf3eb29
8DtdT/Vrxtn2upPuv7qaN8FEIb11kwZaCdNpQTmCbdcB6YPGkdxbP1Ex4GBlI59/px1i732FewA+
j7varwEnZgkEM9m0VENDtxUxoKU6NizEbRoN+2uz0ir0xf/l35hMHUyljERTIihFBkE6wk+AhqUc
VPWS8qV2+jyj+t1qymFhQzY4cEHw3UyDzhQaeE12oGS3PGGnTUZ9IPd2x9CCu68CF9Vr8OY49prm
9TC/MGnrRA9YtFLc+HPhzXuTIuMNdn8G8Ei7po/0W7J2kz95D95Wz+7CQXjeRQyzO6R4jmhYg9zU
IymOR24lmAspm01Y4Atz9SE7FNv+78ZPixysQNSU1TN58uPy0AGel+Hh3W2CTS6Nr30OEQKqla3X
me/4P+kBvX8Ey9jQd0DaeGdy0cly/jeyvRUnhx+xqU7z+q1puB11I6t3PBoamFkmVihMRKtDHqPM
BBPqR4dHwnDO1jmZWha59SSMuraEAnwTawEv3XXhh2o1D1BSJt47mOK+Ty069t6QbzXWgFyfmXC4
CQv2+GPGep7DZ5BKDpDIjQqK8/oiDqcfnsfu/sRwvQPb97luR+WXxX9OR1U/YPII9jLa/OkHiK7V
y4VzLIvNe9g4VFluPAqbFLB6cn0obr+sEY7hZOUF3GkGerpqnYxUqimhg+kksa+7g11DoxGJi+f2
5Q7k4hZ/6uikx0e05iutmb6Uh3Xu6B2Py1BO4PfL0vPTKfMRiB4QZTsEE5U21Oyc7zJFtiD1Nben
h5iDqt+J0bmXWQVJ+zfkB43yrOndim6RFDurtYaPmNOkNQSoTiX75nbNeUXrJ9rkSR+1WqtQf/NY
PEk8rBFaPcdAVdyDUF5cXClRjMb+5yf25Aab8XHzCOE5qI4qREG9aGCpSq+xGNcpGvkLiX0vuC1T
gzy8s6WPAohUZDd2MGlyvrW2jaPSj8vzXb+VG6jL7Xlqo1g+LA42FhQYulkSvKRoilVmcCENXeCd
oCSlepD49k7APtZu3rHt408WJZq5FLy34OZO0dOJQ/pA6RQVEj04Kdrsnce5ZCV1bkldBgl5AQxu
17str+97O4/rmhKdyDnds0q1VpRIc/36NUcnygQGdxsO5/xk+B13mEPxu6NWRd4qyA497XIdIPAV
oxrbZ0HzPEHOD4AkVmvZuj9YnWVo3EJjmDJzHDYGK+ikI/WgusQdhAjkYlHrkUfN2gi9WV7AV5ZO
3BRB86w7tq3Cyet4ewJKX+7t2VLyxHQgvSRyRD4aBq+C2j8KukAGCdGLlVo/oi3i8l9nyDQTBqxL
o9cQ49CzmP+xQxnqGeOHDl2BM0S5evX7Y8lxVd89rwKUlowJWQFb7Lo4685oUIco34bHT7Fe3eCa
iHWt7va3s71+H3wosip9a0xILztrNoRn54xQ6TFMi407rYE1GOCh6V6yyazzjcd7WOWSJqMQpMws
v5JF9fmh1W+gtCnZMkxftF5vjq5VUjueZHElnCx8ko50r0z171406uf+8NGrOiNmNQGe0SW0s4MA
P/1s8VfxYNQew44eccIZubM+v3eepwebZLRXQK/c4ZHUA2LrWpiggtjWjP++hSAjq0Gk2g+1Wqo8
Puf7pAfCH/cWzpWoOQsqQpKNRN5Vj1a/199lB6sjdzvVYgPrWUu3c1K870EqAhN9Qa3kQ+tdYNX6
IXgC0bd5hJ32sva+WTL+qDyiS2CJR9f5sPx4lkvU7dZa0OSIH/efySmy9B29oy4jZDkMzlNmXurv
mRlAxlaK9AdYTUxMExuMsvSRDRx1tLlYl1i1VvHYjzveT08XDYvbaYgA6BtzxdrFo9TgVZrNLSZy
od0vWk4gd1ooFOow6qHLWH7LgvbRHGI+sl+NkYTvR8enWTQuAGQFBBNn4J/qf+K2vovR5Q5ZcPXV
kJLtUPA45m5J/GiK/3+w49zTgxmBsWh/aWzvgA2Y3Ygf3W8hSAotKQ4VR/Kr6MxzR6nDIp6jj4Ct
XdMP4tmLufU+mfNil34hSzhxUWRVLbL5K7Dz+TnAGPIpA02wVhHCbo8kxvoa4iUwW7yM2OpZDJ/G
8HKQZLL5f6BvhP9padacZSKYjHzg5Lg1WTvoEXA9R5vidScqAN7dVYrMsjHZrS5Uc5+bjZg+NlG7
62zV3BP3u/tMsyN7YJnwvb8tCxEGS22IP61qdbYPWCyQ+AC7soM/YbTlXdfn2ktPX4FK/n3QvDKF
olidfpOufO43GksClLTfuvbAC7oO+nvWtHI4DzkQq/CPnBtMboT7fzKXUIr0U3JW8FJnifE8S/1t
Ewqd1gdRzsIiKh4jQFzTth+Gx1R0P4+65E/BkzxpSOkx6Z559ep1PpN2hIy06XpU+qJKJG23akbq
ETOJFMR8PCKrGx7+T+rF2eFVUC47gdfCmtp3Jd3+SSrwT16k6Z1cBeuF6uHdYxj6jtvdaYV23p3b
ul496gp4XXPZBnBzjXHwUoR7IfsyGoaO9irV9knlwhmuYtaU0OO8VzqCNaAlziWCsrSSZPJQYq0Y
Dv0L2oBR5hxMeYaHIeI7m26GenHlXl6YSJWUAp1kQTd7pdIQ+A01skm2/sld8iZjqrW/7MPTz6Rl
F0GW/HpzjB+aPyqfn9OLhqUeI1xqfNjRTqbZBljgqrTBF3ASxtYksXKKgoaYYe8rh8uMXHkKFPks
ratu9OhRyRLLSXqiCWHiXef+JOjQjM+GFsmE1Dya08k7n3vt1HijlFzQd6nTRwxU3B01ewHV5d+t
hDAVNTPnsIvA49Mxdo4mlqtPCkDmtOz+B65G7inQtA6gDsGGAkRLQp0zE+4ROVsIsClInfyt7F0H
XSF7SYOynU+YacAR54z7og8RXq1wZGxHkuBr0BIJXtbFkD6AmUFQnd3MlYxyqUImywBSlTvCS4nV
c1hT621bUSqHIXf1V1rDGMYUHOaHDlO2Vhh1uEsy6LUYBC3hUrbpSIKETKqYUz8cH9xOklti2gPw
Uyn5oJyNLNAhn4lq61BVSGsZyyrsZYlix3F2gt5dtjDJwai8lE2Y5MPJcsoeQlsKrZGQ42hMTTvd
fWvkDGxhD2oKe20SiFU8RKs1ypH+FzVgY639D4jVMfTP1Fnl/TzgNGPeygrQyD3OGlD5R10Vifvj
0eubZitCeQZb5gnnrpIS879qzbEMMNf/SmgEvYGWiB0fA2AjX3xzgWEZwvhv8kAsUyCiDgrmBvBh
argv0dkqlxAEbgdc7BxMPXX/OyGv7ky0j7SBEEpU9clXT9+j3VaCd0KJDWnDanj1fhUUSQtnYU1c
Obz9Ep3Z0l+2iZ21E+H4qyk7yRD84OU3sPqzK/cyAw/x61ux+15ti6x9bQVDtgpBehn6PhKlXFAg
PUSvnZzGwJUgK/0SIkc9uNcfiYU/dZwQEC3D5nsq7ZLbx382RHbhssMRhPMUnotWq6oDtYk90svU
3mzNQ1gX/BiUjuyH4gQRRIFNDXXwRnUhMBNUsi1hHnDtdyR/sLUBuCjbD176JyRPhMExpO1FSWkg
a75M1oVKL+jW22Ac5nPCF/2LL/Ygx5hY5CbFyAe5JAQZ5mwgfkAXKrPZgmWqkMB5iI0jyFIYCdDT
KjpV5yW/nnlvFkuQ6s5L+8w08/PpXBqVEBcC4aVRG+Q7pnZSKVHMqjneJnzn09PUu2O4nWPiQWBj
jf+juFF15bcv4wfZk9kBEOj73LcC+XUYwCSHR909caiZXvooiAZtIjZ1xM2jPLtxjbI17EF8KMvX
6CN/MvjHzHVf3TK2UE2gpEvr8PT7VNS/RAL1svcV5XQIIDJu8FUAEBbN6TiX65fCB8zx0zUmkgK7
kvHlh4iQlcv5Y/qgBkQ2Fj8BW1XIuOyzADbN5VLANu23Nnv49APuHh+b4FDFOP1guM01KQjptP3R
Ha8Rg7EKWREZmEObC0iYUEI7UOjw8VcsGkiygv4ICfBMm5QhcZeUe59QA9a3HmucBzewSWZPVPwu
ZZocwleAG1VAR1VBxX0MRbjBDW4EPoZ47rMxqKsIZRd5Ko7jGyRbliC6mu0rxbgtNmhr1COVDYXk
RUzxCD0gov0ohOIkMqHnbPQbXfRjflA+NkF/es8YhO0DineSM9+H5cOBVIn2kmIdEWf3IpVrkZYd
Q/HJV48ijs9A1G0b0cEplPJGZ6XvYdp4RK2rXljzBP8CPhSQpU6KmDOn36Aa1SP3xBj/F3yx41Ls
b4WYa8GltF1ZfvPp1L2LubS8FsuctGpzp+2pFLtgByGEOqlSoNKJYB8hE9NIxD8lG+F9ZB3jTRm9
oVHR+/aRktwD6ABdeZf3EI6WWl/WRIJM+awR8b9yqrETqxFb9DJrYqrP5KTb3VZokNr2L9M913X/
lYBqWzNlS6as3enqsWJr/F9nNPq6MBy+DHyF7re5uUf920X8lJsNiTCZBKwHFspk4Q7mkdZK3t01
fSlXQ1CPTCbJB938SgJre6KHDJ45T/RE4yexJCfKR2uROmy+6Wykc6WdfjJbUw8aaNGD+BrwGqYS
ktWhyHd545+8b8eONyTvjohG1n6alxCXq6mcPkubdJpUcIma0xpi5JuGM1N/UVQsDIIqmMDnjXU+
yc2/Q8bH35CpPs24wPpX9k8kNaRsBsYR3np6gT1VrBEXEZdgtjMOn6LgjqQl1UETrNEGVQ+RcBjK
PuVqPqpOAWtwyk6x1rJlmMysry0R7pVGYcSKwef8yccJPmoLTld+q41YE4eutRh2BQzn49zSuUmP
p+1vntbrKI4gFakGHYMnd9haJ4r3Grw9I9oK/0uuxU+raNmeHCF1V8pariVZh1tR3slYRbtEkv8L
oljQbmcNmraf/ezelbMFKg1YVTaBuVjSuxdg+uEyl3/SO9vc33ACVXe6F/wtoLbKweBQzpcsbLYE
0sjaY41cZRnEW65QxDSxw8E4Tf0t3SHtZm8wmzSmN0Fw5cQfqzHS5hveEhgfbyKORO95nnlxRECe
aoIIZHof1oe7dAU3wS3Tgehcfj9ThRAahlRNTaYdm/6WFMz54un/tPb2Wx9tlsvtchfCyTsbrlnR
ZFXE+i9qXCnmh0OPol5V08zg17QAr5fuYA8uN6jr168OzdQ334BFgPDzdLusvQqweVFc2DGBeLXn
gpMjnwyg0IVeoMerXtdibf0RNv/k7r82j9/5tj00fsVZ1PBbJUN7XGxeSbbaMXaAcSeae4OEqNyE
baXQIIDqREPX+1CoajFXJGQRK2oRn+QRauWfB88ajJ5S8lO/LAnQTOU5aQb3KyMWmvWg69TK/T5i
0xAZpNjPoA3cvM2wB0R/yR+c1A4lEuYekTB0VgMsCtEeGLozIXBnkFZ9IjVWMGLdCav9HU8eiZGt
cY0QPam3fG56QKZ/Jjo5GLvRFiqRpo/gG7DQgKuT/JSstNhJKXlFLhDnlPw3z5zRjR1JFA/PG6tV
+6iNchNPpT0Tlq46QGbnB/Z0LLXoVVm5XYIFDWuSJKAyszeYKhHfVD2R7hFRMA8saXVGBZCC3qWj
eijvqQQ7S9DfpclqAsxYSw7H0AxOZNw0Sl2KbZfxxvKIqvR2opaghrCM9OaVuvSOppOldWBqAXdQ
A94bNPBPp/7kjq0h6MkS3CLMM/8V+T4fb6g2VOdefAGx3wxCNXjKry7yGH0jsVR8f4P9GBIg2Y5V
mgbi0quxIz4qd0ts0TtN2Wqv4SL4e1xltnM6SGDRXtisuS5Kv41/Ery+oPOXmFaVeHDeW/HtaJs0
AR/ApQqmdt5rqdwTg0oWtouQKINz1Pg1gcvIg14WBdog3/hPwTiJ5DMfQQIXKpGrQ07jHsqReDRh
2bj8lA8s1vg3qg0DIIFVNtgAMkf7kp+Ro6uwKesDA+i2yHrJWhBMsOtI3SX3WF5OJf08hLoXfeCf
mD/JYNMFaTg32BlREE/yeTBFzJMR9N10nkXR8UiBy6CY0oKrK4PlCuKNkhLEW2ZkImZ/qZutRMyW
uOz6xlDCzSsD0/YUpoMoextezrTIJOsvJXRR/bBeMdr0otFML67WSbLDpfDoXkiNyePP97lUpJZD
sosMDJPx4xuUglt4ekZDY1Y9eKcCERX3uzGun1VWzLPTe2xjaPMFmoeMULqjujZMU3Me2qUiM3FF
1jaxWRAdlbtWErGFU2IIhguvARQjREGxcDwCrNq9rDGeDau5w3t23sHzOdy0LEbv1fZe6pjlJLTy
Co2oYkfgxNfKCROmPk6WlJgRjsYtakwGMIQsr2tNrAjeNE/bSBPW3GDzUjm7AvdCmOvTpiTQzArY
ephmt0MjeyWwjlf/2QBwEYDeyjWrqp3e93Fz8SddPNeX+hKOsCPmpGCpdenomQig+cr/OCZWe7eb
VUku2fkwJ5CPOyoSTDq21rU45M4kvyCrqa71f7rr6tHEimAJ5KZUQUs2kRBUvubucSmmhAp7gt05
/5s/JWnBbPbTiPT/jD09Rgze7iV5/5u9tnU3rHklMdKmGujcCHUlrajbOnfkm/L87HyieGsrYJyI
lWIPpPf379iAgBS7I5Z/Ox6nOz5uZYcFClvT48hkPbDZwtOHW56v2qpDDlNiR1fpXB6uZ6P9JiJt
1oZcGzytSsYTMnn9HwIfy3GoIj1E5Tcvg4lwikCBc4oPxwVPGd32IzVvqzBsaOB04SxlPIpNbrxy
ZODyqYiCD0c5JTr8muV60ha3OGaMRD+zsUsWQ1Zn0hTxJl++dAvPM5xmn/9DZxgbYi6sChNRNTb5
RAIw/Bqw5uSj9gwb315JDPHSUR7xEl9C4hgy7AYxoLwWSy+arkapFn74/uKg79oz40tg3xyNSKBB
/ZzurhLytPBhc96FtRhzXZZpv+soBcfbPRw6HfpwphJJGUN0RH1Lvbtk+v4rftijuQXpJj/nQGju
EsklrOzMUCh8xBoiR4Fy03TIXUUOjx6zmkxN0ha9Cc9Nla0fm29NnEVV05lRQeBA9M09/cfOauNI
k8t7O7EoPXQgSGfNDtTgcmHpocHV4ihcaNmvPjgAbPK4OuCUm8O6XPr6s3HtaIRfvXRsH10ccuDA
2hlm4jPwfFowfjbKqEWLC3p7mlOZ3PU3hTqMpz1u6WP9Ir95S46zSgyANPIcxV3IP/qqsmJzQ2/m
w9FquwZcSU+Q0UU4nwPpWx69b+7ZjAI5XzCbxVsv+nMzX4MY9Z5cN/YnS8qEoMlCkv7poyfcwnNL
QXJkBgAUnt6grL21w9+b0awjBv2LaY+fkQ8Yz+GnVAOpCp7wOLI6R7qjPnY56Ydc9opk2V3BL0Ig
vZNStVTloj5WV8lzqMura9hnwEy6ocTAigk7kH7VHmktPZQLLFJK9nIa20e9wN+F11jV7zG5j3fp
DsRAQ/RilCT4SXhnSgmFJSYmjxGJaHKSd9FJ151y8Wt1tWDoI7p1KUpS2vIEPVCNBBuXCGcSRrfp
ccghaK2RsRvlEKDRvwVZ9AUXW9JpECsXeJedbJhf6lpTGGPqz4eGDInL2j60/6cGFpm2qAIZHbvx
iDusA4A4RSat5Q4oPz6nf4QSUYjcrNo4aqZT21SiyEYbWpamjjxtovuPm3db2Dw85q8cDMKAisTi
v0/qX1T7sbGEffdYgkpvogtZMHT9KOZZPJH0CJ+ZXmbMayI0ElQw128hBWyw/eCDbd/F00X9qS3f
2t2tshBy703Q6/PRPDYWw8rYd/S+bn62fDiHPa3YfPn9rohNGJsrpJbqPl9qRiI/g7hRSkNtUwi4
jEAhcbOk9QUHMYY+VXVOKfh7Uf/e6CdG0LtX04khyoACeoPMjfFmZ0HjYIoe/11jdS1heXGsGl2e
e37ZApX1/XQCIldNTAyNNdNBpRlZaGGw13SnAFwYsohbFsU74kenmUaC76TiYyydXyA0fsqdS89v
SpsT8BQKZ8b+InIrPlV1AA1doKtuRvRgMOoobDummT8mO7X6s+KTDgKvCECPIOQQeFa0//cUMSuh
hQzSzViyF3YUFQD8YFEGvJ4O4v3ihwb1lnqhDgO+GWxNGcBEOkoQAL3asabY8fsCACdvmEIpSZ9r
Sk6bTXNtpIqJzLl1V/d0IueBbfTioA/ge4ROYKUxJ0EQ1WjDruaLb6pOHnDAv0YKyNbnEHp9Jp14
+DqpaNy2HESI0EuyeZBWFuIQ1b5LRNJKYXLU0eEte2LyXkJpXykJTGNjZ6SJ6LOSNs48kaxZpmWS
W1+KCrJ9Wj00PTUTJRxU/iu1/E3zKDc/mqTeAaR4a5nk5Nl1crUdV2qTwvF9gtV0tQW7leyofh5I
tgKqq6efPsiy/LTkpsA06tA7Fj8/pXtFxb2hStW6CO2tVt7Lf1G3lqIbKAX755mm86DE3x+JpGYn
wu0Sk3c5lfyCqB8BqTPSDZ3Pep24++uvmUvlUMPQmO1NOS4qj3TL5gAyOWSzP71GlfCh8qysWZ/r
C9syPW6CULRqpMUkWtd7IP5WafeYDG9f5DNrl/mwaUyVbnHrxqELT3i8ebvdHyORE/vYxtznOQUC
/vnsFfQZb7aU8wS+r5K5WP8jvmVcEp0vFuDpWhYqiS2G6FyHw74WqhWSAY4JfUuQrxdDiV/NaHlk
hn3MjrwtRjfxkEhEABWgzADWhrikdnLcJcHs96qxsLaSWVmFVhFyhIpGhTyQ2OQnTIvvzQkgQh0Q
TEFKj5rPMHr5XTjYryb2lN0wAdu4R934hDKWExDByqptQksp0aVTcBiCAsrfi+lc/dZCI7qiw6jX
My42oKT1n1zjr5UQQzhthShfzw4fbdsNEwtzG7U61vFkk5rctRBwA9LTy3HK1EBVP1V50nQTCN4/
O5AfMqj+OoWFClOPq8OG+FieupbLFFxo87wRbKrnVXE/wVMzCtnymdYSjB9ZvRTLo5XHOjcpAxzW
qaZMrfFO92AgRD7Ci+vrHYw+WJaVKF3oz2LXvx0uYgBD21cONaMTuEoi/T2W+m+PTB0mKeZo2sAw
SWvPimP5EA0QaI1wbAqxjxJStYEflzT8nbh8H67zsbv1YVMxhtPV8T2d5VBSA0mXW6OwE3MYLmKc
XyMUIgwlDMGNLTALrkPCSXpCBbTnOmRcx5cn7ux3DkMtyYUtbI+WcNT7uCbPZYFlkjbPTVebnODk
j/omvd8eU0IWNgjIThA3OwJq9O6ZXDkAhMEUhmLUQ9VUJJYjLcJs+Gy1/vViAAUo7UVutCNwsXc6
HHJCY9SgK7sEWCmCOirf4/eOnIqtP9V9dpjEqmdSJakYBrIdeBpk1niuvjIKV0Rv8MG4S5vR4Kuw
qTSYiLAggbTwBrnkgljygRBfcdJ1yoh6B3tUOIHM2tcFzAhKDp5PpPbPipjY2VCZUyBABlrYNDM2
lSimfN1yE/U8AHm17SVtNoBYWRSYAbtNbS0FIu1MlqxYv0FYjjqA3Gd5s1panQxhINHu/JSyIv5I
FbiWVTeRZTqU63v+F58k+I7m7hOq5ZMjulV2wVAkLkn1eZnQ6HrY9HkcG5zxLEZNd38XatKzU2N+
e7FiB+Ob9JCF+7PpJfUy6b+hvTr3MvER/Ysl/MzKFZElUGz7XSF5/N/V20Gu5YVqjQuCCIsHFaNK
nMq4lFD/3TFWQgXmOQFMyxkaKzpFzX0l7COh1cYp10CaPmDjaqC5iVok5cOxK/grV+UdBruA275r
VK6jl77EIp+vRwQ9jUyEJYp5NqeKw/WsYDwk6ZxJMcQXNm7Mpmpnvn/9tj2RR84i9nW/Ljt3j89q
SnyPKB20wJmNTZmihFq2i6jIFQVlYOylP4sOr87mTiZPfsBOv6lUMyLG6D4/sNYYcGaZmtNwHDwn
zadqkVig9hHJJdGRE+8L/9dT7R8FcnQZimlGQYBeVX1FB5/W08QJnrSkALwRNYKfMrGHNQnAxI6l
LjxssWv7casy7QjKVSqD4O9VkY5dw9csQEp53s63q1EC37tL5rTmiwwQZCMsPxZWk8m8zvLCgH6Y
t6sWb8MW3fDcatrhAAQDEHbGEhAXDyCwck+9OaIn2B6PVZLJ+JClXlxpproyvGiJsd/JyC4HPYoM
JKGzG94+bRz1u/0d21QHbZ5JJfb8U1QmnDjVs1cF9fJeQ1NShUibzwNrY3dUOImFnq62Ga1H0MnG
G0hvu/onp1pZnvkQ0c/b8/Fi+gQHTftm69xffaWKtZgZTNc9WKioGuT2RLjO0a2VBa7Pz9A+MK+R
NgZeLsks3uyQabu4UeCKI2JexymMKzkrDalAvQuHNfut1IF8KSKzbQ6Taa2Gx/Vre6bM860kAbwk
sUhwIub2oCnyQC4SdCQXGvJew39ZYMri+dV+RVJC8sB9q7nSjlMndrZa+rZ1beMq9ulkLa/ucA6h
icWshQe0xH8NgD6Upue8iPdrE0McP93xp0T0H15XS6zB+NZHH75kz++EBqwu+XEhPTfEK8zXYbuQ
hOVtDZO1WUAkrnzQoJCCFbrgYKI65a/3hGn8scpx2eLpa90VqMV/lX/5Hc+DJPmpX9Ud4ww6Q5Zq
E2PtQ6sLqbbpg0XMmtSAZQ9kB/ZyfGakRg1v2ejy0ciVH0E204FHhx+M1FqTnGtOgpztXLtABkco
1rHApUwom6bsEd/Ktt/zgpGg+4YS0mCx23vlLdGSSLHLQorVffeYAOM03WsGTdQmfkPkHJNXCaeH
bj+mTtE94iumsVe8kgySDqY+7hpDnEKOzRJE+gpOf22856gfKNbe6cF7qnpx6th1QqBY053Qese+
CI7QM9Ap07CWzykjya10G0WQ3k0t73a5Pp3LetnnvcH6dFTEWbJmZcEfmRLqeFbzNx2LBGvvkP9J
OQvBWAbz6rXmpGi+nyiDo3DQJqcMnfcDDDEvByr/iTS2VgJZobkcX5y+cdsoapwKC8aSGBdrGI41
74/YPowbEwkebT3SPB9dMdgSIlx1VwS2W9VN0HaVLpjuH+BhlMKq2skiuugIzjMlieQDVOapXZNz
ZtAHwHCIsQ0SroEbcKjlQBhE8Sb6P56fkghp6mD/846EGr7O+o4HaCGs3kC9p318z4sUaCm5jBnn
nsFx4obdNF7q7GXG4EH/xUr+rBFU53UuqRTu93M5xovUUsErqD42RXJwM2T0dLym4xaXFgy+jMp7
OedMBiRJmsp9Jt4DXB24Q3ZQJLM1Yps6n0pWG+NIBlC6G+uMvGJ8V0WDv7jmLfzYGax0Wj/BRR4q
XITdvmuQN54VmBgztsydoXrAAGvKWEB5ExFHO1mzVYivBo1m/DxGMsqVvSIuj9jYvY57uBTH8/2y
GNLymjYv5GwG/8Z6nR4lfplW3yPjkbN8prPSG+/qy7UBKd7AmRjQ0UBw6BXfNPJeURJW7Ru//HXC
UMHPzKkpwLzbImr5RIDSz4Xquu03yXWmYzWRgg+gpaS0tsEJpJAFWLgLzDb/CrocSPg4RDXZg7nF
ugPldM3RoXCsBKMy92KBZijWkaHDj9CHcFWOo8s3IYJePBYIx34fxD3asvS+t580q3qykhsHRQjm
dwBR4LGZDIxKg7QQ8pKvsNrKNMT6CdrQlgY4y2QhKZhJ9EGIcLMYBNVncNvPDg6Pl92St9OpBYke
GQ4P9SQJqB2nmDXh1TqsA4hr7MPwd+KgNL9/uUihI3S8QC/YTNVcC59qKTNvJg3nsLOWhMnHuadj
viSRNLWPV/N5hYPclNUvstjQXBZH2sCtIfH/kHvANY7yin0Ugn7Po1EFjQSQZ87RDX2ppQqk9jul
QND5pYqoWs9KSkWoP61b6Po7ZlL5oQMoxnw/qENS6EMhzeDYf45cKYlq0ADewCjV1Rc5qTnO7aOD
17G+WWY5E+zzLb3x0fFEQyUWxs85OSW41g066xwge3VsqItIVHC4jBG9KDUNQ3JiCteEGBT2H6h+
Xajzla/SoW4TdutBhueMzxgwDZmUakhZPOpY/eeyarEzng+1eyz4GJi+yol/Zluw1FpeHVIAkkwQ
gaqfPh9/kojGf5zU67HLLw6+7M2gYge2qFTYlQeqvwkWCK4bnaGh4nPE+LyW4pj0J1wKq4xt9eTw
FYnS1Lg+Z6V5JWnVK2ufOWyCKSy2W19TciZCLqedvDfLDRx61YicXScVPFAgG3rBS8MqFCATgXhc
fPctbS8lkxwjC87u8Wc5utx2KO5PiFqysIVqmFWeVsjTxpM2LlZ/lF8LeMQn+74+TaL3HgmMtn/h
mlK5BUWsoSlNutLqQaKfcv4eXI+N2PpUz3eeskzXcmaOSc6cOuMfMAHjiCXveQDey7t6N4Pm7mG4
xz4c6G27PnMiKTjiZ1Ir54+5gI1jlpVFuSktCsN/NXvwzAGZmArFl00BjUqt+KCPx0d0azTichwg
g2mGvQoLRGyddxiIjtu28SaXmd/irRB+btdX8W1ckGlwXYL0cARfN952sd2DYdXgQ9TAPWLQWou9
iwaRT/jGDKf52ypHmrLx56Xhdz16/L1gL3Ehn62yxIJKmqsDr7Vbuf3SAdLYUPPWDmGPzO4/x1Wy
YNcE5RAff7NPMRtVU+4/xxXk9JvTQgF4XhzkTQSb+HreiuO90iqVrxi5vWmr6Zt5AMkFsu3J8x6O
1nPM97Ge+ynYRBaG5JVl7XTMRjgJA+xMZ38qiAQY5Kwt/SgxaK8aU+k006fOsIbvxm6PIOegbrHT
S+uSSqYRaoQxKbMCd7XieKByrnuArOfZZY96OO6fAtFyGm4s17PvLhSY3n5a2v9klOX/MaxOK9uq
3B42mH0YR9rFSrfAxjcTdEr+r+B7fXrDnIQkOtxG936s293veYEBc+R59QkdRR1yNpVFtdS5W0Yg
e7OhEB2+Sw8nHXMewmA6AZNs2QFFpsoufY6ZM5A7NorpRtecU86jRJ+Kf0OV0dJaX1vF5Cq1nUXC
xa3tua6y4GsBvfAE29A47vLvmxNqRJkqkcOWGUhoa1Hp2qyjX4ZRgnmCHNI7IKQVKNdVEtCwpVEI
EWpQyCLKDxdxzK3Vxb2tO4Dv3SJxweqyBK6C6AnyGrP1fRwJIlzRgg3R/bXfG/OEHrapjJtf16hz
l08qLPguvEdTUpTTYQctnswvuOWjRX/nr2gLXbbbZgsMmSlMRUPsG5UthmwYw5n9OIBL7I3yPZnP
zHJ/IS7rIF/JSbiAUqy8P6/aRcLH+OAuC+neC0LRMLX6BfYZgZFft+BETnQtCNTSBQkkTMa9kJ6u
RFUUsDx6h01/86OapDeo9JOFVrbFz+tOt9h4351zKVk740WBO/6tuHWPt8Tmcfa56d9i96BzZta3
tzrNh9nTDnCsRAGv1JwtmNp9uNC4aMy/yXow2EqS6vg1i3humHZFNHbLdCn+DSkyYsytWeiB+4D4
xmFxJGVFsUmDWd8Yixo/O0jsONQG4Tzgh/YmifFQEiv8MB77Q2CZx1Tdz2E0gr9Z+Xt9v57zP3HY
cWRj6b679LiXseT1LRemc64mgjbym9Gx4SRx86tMr4F3g0X04s44dvL9JtStN8xT9guJYyy3sFbh
mCmyX+8yJnf6biYa6hn8NxctLmoCmKuK1I+dLnQBsIROpnPrtnYUNQYhoUwAtlX1tuQEfrkORDnB
mY6BH232yLeQtPalfmhZn8nsn1jFWsHBc8Jh9aiRafZVUEOHZ0mbAJWtHRkp2pA4h0sUtSjSHnGS
VOg16iepUQr1dAb6e9dCttd4r0ZfnYD+GPU/SlysP+JRN5TfuTChCIuOdsqVfDHpZ9oXFscJYBu5
pI3tzWBSSdTOZiovm6evGm32fuvCgcVM4fnzxw41i9JFFRdL0VIGiWnSewpxe2dFQ1DZSt5r0SBg
xPPNkZdp9z3g8GLnksk1kGWEVLXz3pS1DVz0QO2vrEOn5ncMBYZG1GttyX6U8LmDxwar2nl0MjF+
OQ6SJFpPTootIaq/TxUwE59UbFejw04BwDR+tIw8xnQLMVDz/w/myJRf9OJyv+jzUFnUSDh/sKfk
T6Ve3tW36pFeqCl4hpUvGWuFnj8L9xIIIIoeGt2NWT2DSwb4mGd3c8xsLyAXSrGhRVLZkCxNKIov
HEjakj6f9216VbQd0nRfxNAE8gJiTp0cEsXhtWoehlw1d7Sv9zkfSPIgFulX6a2V2roHc2Trc0qR
5ElYIvieF/PlLPF4AyWUSqVg5VVXv54jJV7ZFdnzpJXpmQDCxSnsONKAaApfwpgC7rM49gY597BA
f/dLac4LwrEqVWD63Q/VwONPvLp54f7qXgETHpT7tNF6EXXnCWs4wfJOpTzvhPow8pAdmeTkaL1Y
jqi3LCOEyQTmuWH2kLSmZLdIjYnPQGAU/EXbIyHXAe0MOGMrxNcurLItQ2fcqfKXbOuzvsVCCtNN
Z0vD5KKhNYKz8eZbiURnExPtx5Cx2MeuH0i4jducgLWn2W7Jp7+dgg8cNlFzRSAT5IoKmu0eb+z4
pPnW0fs4ysRAasums0oFDRvwVGWuergJcMApZ7XC/Hz1D5WF2LsKJR8DOdzwUrhS3y/Sk5TjOvvQ
AVHBNkCaE3ccC3dKiFZcNjpYMI84cVX9K58iyVaUZVTnscZyoxTXNCQpvauRNbbS9OtxyDO9xZKM
A3MdXiVJW9dZR/77YFEST5+76Tn5E//k0Z7SsfvFzEkqLTyi5n8IdLcxQN/7J9LKTe2hJxuWyrCv
xwxr0O7xg36L8oleeHUPwBZBWb9wJaWpL5vPhtm06//CtbNkdnFZMy7y+TX4ZZ8N9PmL2Pvohb16
VrVN5yo7iOW700+/lb4KXDUaZNrypH3nY1D6t/297+Od2DeCnrn3+XCBdj09XcA0Ui8SGmaGRf2K
J5KHQo7BBAtLLhWWd9q45iJ7qDH6z6GjYQHkmKv2S/yJZlejDZ5cyEpJrcCMXIEknvpN4d2iLmuv
whM3BCStJw1u4ANmu+7wILq+XQbefQ2n/PPUNNHFCLuAurF2DcYBAmxJzcfItDhFBHW2j4O3MEqE
Q8wVU95rJl6fiGGW4L0NB9LZbsm/TV++JPbVfK4ShQ36h3YxYG7FNHYfJ5yN6pWJdL//XM4PH35u
PfIAkW0DflVAQYRw3hnAqErS9sqKZ0g3ZV1vejqpf/2ldMUByY/hZMfpHMEUs+q225TNKoEFCHy1
EagjUf9woKAjIKsR8VRg78+8D/Lyk0KxhUN6zpj1xCdP0RnqrSAZd7BWGbGyoRdLSuV3yAJmsqzl
giJ8RHkub5ylyw3fOpxW3jLAtAKziaKm3BfCuy3yPXXEd+eTgWPrE7QdyJaNNiOhprH+JYpZGieG
k4cjIyVDDwuwVn1MmBve/a08yq7ro5xRiVSqMN60jKxAFpUyYdbQMRNGbLcVMNuzQQm+9H4QbmXz
Ed6L09CJy+Yb3iqULeDCSkKdR3CdG49O7WjSZvZuXv0zGlq9WTwvO36jA2QyIkY598f1HIZSkk2E
kAGwFQAVyl5oXkAlCmTpf4VV+t3zrS91UK0txwGyQ0uyPiYK8Qi/Jr+E8Gj/4cOuVdD9CgAzJFNG
0L/GWA+GHtxmHSYEpeS858ZYjxOJLiOXv/PqCCYVWge8K5RwVYNofSu6tbH+KPZBunjl7fqnr2bl
01PspXGLuB9cSs+k/7rfj2Wnlmzz0pZoS6+yybLvIPzd21t3+veipQXqSspZzYtihVT53p4Yvijo
Zr0FclH3E0p0bLjyNainexH2WgExXDLyxYAYsiXkQgKKCyG4M3YZ7cCy/DGWAZDmsT2an8lWFL6c
B32JNnJsiUiSJmlOczJ1Bf32T4Qy1OKWLYWS0rrCzRhHYUDCoxuf+HK3auqa4wDz+X8FV4dIV/OU
N8ltt/G3Jo0Evq+NESyd9piaBDZF1EZONPk6kHiJGw8Da6pfUNuQ9l6+beyA99LDw25Ay3qkIh8p
ZY7TliTEpBfxZ5zEN+ct9psM8KerXLZXIqEEBNFVoXWnIke1+VdP41JkacpSSlT3HCyQqo38kAJ5
lnykss/MgkcdsBamj9medTG9g8PY3bN6LVlYwQoouWOBKjBRE8dnuklqrguK6RqyqesER1Hx4aoj
elyXQ3ZzsetdI00tpsoHBq6GZwRa949Up023UqxSAsaTMBx0VJkoFDtIXAIHt4Gtn0loA9eaxAd0
RJF96K1SE45QSGUn/JGz6sTpBEEtEwFzsM7EoLaLeLrp36FVOmwEciZ75XbQvIOrs6TO0LYzMS/L
kx9VmNXWOHtEDQuBl1g9Bk+sJF5DgtFUga0iU2/o+O8kDvRcsgtw0H8nsa9JcXFpEZFu6TJN/iLC
Xn2Yvd/tbb7pz8Bup+ix9nXeh7tpDqmqOXXqpdRMfPPVv16Vs4r7RLBTyASxzvQ+pXjj5y4qT8wv
/8NfHv8HyNmx4ajtl5MiWDPpOQMYGSsRJzAtP/9QGdzu63vVRYipzm0+n8XQwpyC/yQ6vXMeeg7J
OrWyqgMT+6SijfnojHFHM9kNu1jrdVjGvmkUltBfAP90szso67kKVM+0CBgDoHJDhNMgrcD6AB5h
vxWuJjBY4ZCGbak9pPgUrx7zJHz23N4DMmQWv/Ozw6vLCQ0J/9bIcthWvgSU8QeLY3viTT+Gch/4
P+X4q9QwthzTESBuArxYAiEry+d1c5gqlEm5lZWvJjquqLIjWyBIeRrlKpx9MU0ZPWge+AOeE0G4
+kD/Zp8kMNgE/FGMn1y42XO7JaOrJueaWkvv/u9D2Qhc9j2RH/pMSoDmG1lfLYSzqeUdTlGSXqYD
EuP4GvAG8WKAjEb3hhxPkWM/lrpmNfv9EdBqA1H61XzHW4NGSsdOe1X8iArIcbB+CmRq0qnVrfRH
LUfVBoxMaFSB77uSUy3t2Bzx85mAqLKnEU6TkGCtY43+NTuIVOG93j7p/csszcaWc7a8wc/iLRQU
Qol/73enQKODVAq5p3vSTmMxqMJpmRouNb6psyoKLAiDTLor6SF4YJfE8dXTH5lu+yaPJYIKp4ns
uDleV7nq6uQwMgvmOf30FWzBYhkBTHYjsl9wAB1R02lS4wNMEvChRJMFo2WiATEEgEpaQ5a6j08x
V3j4ZcqCdKmgdxxs5VjIRHaTDrD8/mc6fH3k6h05wvghzwSJUVIMPXjlVaJ99+KgfsRPw9yJks8c
WAxAbmxF6yz6qbdO5dnZHUK2cUBy9EqrAZVpJzSdT6MhoEvBL38uCqbn6JHw4c42oXUvA4z2X7e1
eB9PO+VM09YusPAIagU2/3+me9V+EurNa2mSljDubezLK37MUdVzUCq2mqtESZzKmNryd/Mry5Ev
5kTCarLk6S+eyr/1ipOcTN15dBqSd0woawcLM5uy8clcqrB8HVJexhoZOyKWbhUE/glxWEfJiu/D
QnQJkH7PeBUAoRB80NpITSowcA9GlJZD+DHG0VwkVRK6nogA7S5ZGxlSgBbVyCMa6ybIg8CX1IrT
7AjdDNAqfOBagStKqTuNalQkJG3VaeLM0S0pCmXvyaNOyHM7+/lMMErbuQ7FPisZSbTQPksbwD26
B1P7ClM8q9ahSWVpKmRp9hExLk/ejdjLTKthoUP3q7dIz76oVdbZEy8RworWZeCvbQoQv1dOtzEm
egWHu6UuQLV1HdMLnBIeSaWMOlaNmtc6QYieKga7XTzcoWUhDwS8n9KMUMXDApL3/slqsAG9wn/j
8UaYWiJnQf4uT13MN6j8XVp4z6AL4YAsKPwwxa2ZrWQIiXNfkR+X5j8IPJj6xxq338d0z1Yki2UR
RnevUT8F6Fb+s033hDH75EwxD2weOGHJoCFQKiMj8VxXAq9mmdF6OhTrpfYT62D7s3xWCcub1Lvu
zfGOZdHR0yJvDtya6+RHou/QkANxPWKrHkOUjyseyHlbhTo2pdP5QTjPJazyhHklvgMN8Kn95syY
/UAi3zK+52UT8Wzkm7j0RcsfJ70rcgj0XBlS590Rwa3zB6wI70j49uqAhMvkNueTtSKA5B9BBuKX
j1dNvg1G5Vq1hbzGxhGT2zlV8CsUm9VY8JIlzDmGV5NFB1QKBonAMfBoY+aC7MWvV2ip7ldX7VEi
8TkXN3YEbzd+CrYGA6tArK4TWrD8BpoZraiF2fNkLDL1LruaXksQlMamZzoglnGKiNbgAFNnvsy8
ScJecayTTKM01GHF4UraF8k7gzaYJth3PjAbSkKyNKoE6+pUR20xJoTI7q3rBeo60u0ywXegQpIK
/+ysUO4rYdfaMtWK1SfXa/ybYrshvlCVb4oX+z08FImkzzXRV6enQMUaSXbDu2EZuG1BAD+4mEgv
OIj1qXMFnl59pZLvWnQ8rh7JsDtQUZxb4T6ns/ALQrZ9GGxg4l5KVDq8E7nXFicMjDTgTEWiJu4h
WYriNTVkRRHTBPm/P82a3LykbqSnREYj2RHIz8q+xwpHGAXeEzW18eYnHT4sXct1G76UXMCR6Gbb
Vc3npKfFXwWhIkI2Dj/f3VzuZed+Mbh7ZAQV4gbQ97d8I1CgdrgAYN3UGY5mmU7qK/h5fpkrg1KH
HGMbLJeV+8gVB+xaX+Ed5ymIBEEFX3g9e/DpVzOsPcxkvVTJPeLSuZoM28QdmG1B+qyKc9Og7sUg
0zzj/YYpptNKXVOmUKaXGkpLf1tHALUG+HLx/UmkpA9uPLyoK84ZapYJIOTdXg8KYNE6xLljonR+
1NMYkbIfMGW7zaw5xPUZ8umySGmsQFv9SgPtzhsagI6wrI+8NpWbQLUqoKeHkBsnV9HuD8cu0KvI
s3tMt0ebVW1cFkvbwbmP02VSoq7XVyy2Ag/daNQaGmZML4CCCOUSwKKIOWqwtt2LuSbekKQm9ybZ
vUQpoYL3eIeyotvbw2a9RH1rURqVwjKXv7GjQMuKuMhnmon+BnTr5EpS0ULGqUk8xaNbdpbc6IqN
ROgJzqk1DrWyI1SKvrFLnFD1fTh3Ol13SZaN9MrqPcjMhpWmV8zNfdmzoaLrrnvo5joRAgfg0zlN
Btcbzx8X+tLM9TxlZemfBKoVjsHidJ16pEhhX5eVQj37nOU4ZzVAkNgrxBiJb5r1qRuipooBX5Eb
bItoI2CnaumY/d37KhkRarHiMCT0oNe26qBB8gmsdiSu1WlVIMJtPL8wD/wuEGRp8kA7PUa7BSE7
2D+xBOOHkdbuwfTw/n72SBe2F99flY8hSDwWJDm5q/1hNsaI/DiwKAAsmt8H2ec1/RaVbYlmNAr7
IirxHSSUgQhcoh1mpbTpgQjcufQr6KCfIWTDQ8Mvm/RIGa+8s/xvXKP3krXpUd4xL89tdRFX+ilB
nhEKfBxjZdukUahrek5absYPPF10dxk3JcIb/CpXxeOzSYW7lL5TwNOfQsp8jaCzuQYThKOhEPsf
i7bhznIALnhWJ1xXy4JXImDCuxSQwD2C0sYN4MpeS0OGDaCfQCsy1V4CxeulRhf2qP0ZouwnO6vu
w7sOU2rvz50s79cD+LS/PiGsiVN2DZGtyDM8fJmAzuHRJ+e5GU6SxwPqy1SawGZxHgF1iMyxnkpw
8q9sg0qbL6up5DFI9UXBjWTMPzTYLG+4xTgMZ25q7UDcJPKQPwja2UCb5DN8PwDtjvXRfiT1r/UT
jwaP1DgPiQar9UQGnzpUX9ZjOTRBIVwOsO7HW8ik6MJ8EVPPRx1ca9CFRk/gMnUPUy8LywNHpLlI
F1f192OPdMVELf25fqsOKJQbuIgB5ZxThO35EVZWHfVE56NyLzFRC0feI5CBPIqULv7+5WocP1YB
n3f0OioDkrHDf96u33WGTrT+NjnUGoS1lqvira1i3rOUqnSUy4DZ+yWmHgaCYxyPe41wt1BArIct
wOgfw8SMTpGTdsH34ej80jKK1ssonxr5lfT2wTRPlI1S3nBLVFepA8ylOfy9uVeBTxZT3BlxGr42
iw97yctx5vvWFvAquYrwYtmwQsgXOFpemdrLLpmhx9SELrUsEpn9dAhoAC29qr/tHU4FwXQvkziz
/rF5qfc48kfUpnUfOduLHg0rbBMKFYlLZxig79qs+H1/7wbzr53Jb4XbveFXgpNu34Y6O2CvIlOR
M4OKGuCcKxLfpPhvcPf4HSYV/YDupp8IfEbxmpIkYY975IffELGa8VO2dgrekY6NEngwpzkXX2vf
dYtVwe8HOiu6L+9Eubg/ix5Ucl2t9K+3d4ItOzQn2e3GDdDYgN2s6VbZGGySqNvWOv9jLb2lehzZ
weVRgmWNbBzDYRqlDBEGgi+ojPX65hhiDEB75jY5Dh+kzY8pB/xsQ4mWUFjHvHsavf3JDxBqEcSk
avzS5jtoCxe9oEcXfGbH89MBFMNQYZrcQS1ySC7g+VY79KtW8VY2ytFRbPOo/CBxDCgwY6q/WS/P
0GRY0icwZc1vFQGfTf3AJCsRcrZTzRyby9hlarfqwxOrKIL3bT18d2r/I7r/AxDply97hTsHzcND
jMumd0F59/Vqm7zAcGflJev2D7YtMZrdFP20ZK3AkkHnRt1ouS+twZcridnv675TQklxgIb9w+Xr
rpl6ASykiRkYEsoGjI/2Q/1OWcEyE/GKrevs8eH8gkO0SfZprK15sNDqKjloTWOE6xjg/tyAneNf
jzdL7eFxoZVUFaDTKCzmU2SF+CMnKIFH6Yi1+D+OvotZLUxx4goC5BO4CNigHXlkYjXnUJ1P0EI3
afaoMWflwn7qSdGhCaaMc7jmOSRCRFOYotlfZPE/+kTBaHgGdUI4mTEBVBCTrsXImOcniRemG2fg
uXV5PW7QR8WRy86Bzgh73DQt5bxPxsS7ucrV4W6OZDOzFUgrz619+V+pjOoMzV+9fgPerO4rd7FV
DeivT8VISGk+DhXLfGQOdtJVPT10axBhU6dby0BKUNSrH8JRd5O4sJ+TVd0W01kDiXZtv1lpz36E
qPtSpbJ7Z4jJeKpXRTWkT7gR8ECtnYUpceK7AuLG8Wleua1wOtiYbdJpcWWV4yjYITCfuJPCEX4R
MP6XVAJv7eOreyBy08o45nRyFUX6SQ+GZHWbdKCBANOpM+GA/FJuBdsKOlqT9Gj8IQUba4nL6R8v
wUKGGuhqcdAT2AoyyeLqVyo/saof0QcOOxOoIk5T3iejV5Gb7Htvvm4b1REK6Um4XgHAwE8YMTEt
hLGerEDv+zO7Ethz4VRUe0f1Loksz6qY/nF0l4+j7Ge7EgjGrSdoxi5YIgjQhfYFYIXV0hL8YIj9
mggTW9fRUekxMqC1eQNGyUf0qH7dG2DkRZtcpVRU+UNplKWcW8xxidZFPmv0ssfBKqHPKkBTAzCz
tE7OrvAAQ8CAq2p43gUOOZ5YOwQ/2J13vJkojeuKWpdAzAClnsw5c4KcYLxzNvTqVRM76BEO0Hrm
FB4b8Ce0bZ0x2ej5rOTshSzIRjhg4lgJJG/GZwjnr5uODdh5p9VJyvpp/Lxauj+fcIalHWH8OoAO
s2XmlpG64X8P8aj3Cbd7bXCD8dQRq+PRyeYi/N97M8HQYfuRwVnd4L+aQJrUJ4lDe6TYIB3ooA3q
b2VvJkUpOGfmNDrCCpC5/J/B9/L2BCcXHVDfXGWiYwYHBLUVCJwZOda4Ag+SQRRgM+jkZSob5zRh
gRKF0ogjy6PG1zKXJZ9Y64gFOUsmzf1THT1rkGZr3ejTaE18+ajN2rETDQxaVCQ37RIKiz0zrQCj
OW4QGbxsjEVT7RNXRKOEKGdQS948r+PIeXdkCzaA66lDy69wXOQTDvRxu7joKOGQXn4yQHpBQ5QV
9Ma92xIaGy0guvsdrh2OeJca4hDx+TFwCIj1WfVYVtTJckP8OX/ufn7SPXt0ycsBXbGoOn01c/lx
Fp/c1ala5YfSV4jC5PvOLvM4nhqh6eLn5hPjPljmG+yKMah414ihLClJvulh7NDEeJbJqSkoHq7l
AleIo5rwYNPZ1QJwOkZNrQdaUDcFdQy1BWeEb72vJm73yxAPLel36aPyFjW7BkBKahhonkr/HyY6
r7HTrEK0BkwdyKmUg6Vl1zp4JwdOy/c8BTALawhJc2V/T0zZ9IQLQSkXEHDh9Ay8BXh73fo8gvCV
uOqvE5WXZO8mcQoOlKyRNroLauRRLns77NWWgafGWhiYLFyoUM+ZXPHDa+R+Df31qLP1YXzER88x
1qoJ+VmOFuVB1ruQ6IW7nNsUVfGJ5FsfqV020WIRiIrdT8SEr99J1D38pSRp+sgsIK57em+pou4X
AjAzjPd1XehVvffy7hBRT5XQL745Rn//LTVx9L3HyBW9KTg/OfVe3V9ysxyiCWZ0WmvmKfX+86qQ
EW6hPCP+2SaWdn7+coVt40sxr2nOxcwegxiZry86rXG0R9bb+Pk5wVcnaOkJncwpHctho75bCZQB
kyC/wEWZl6KiYJCyHJWLivLXTg4FC611jEuXZ8M9AA7HdbEncB8D+lYVYh9CJBFSdTQIjsayZOoG
IFJWnrCu/L/7Ma8bLFvlNBG+qNQZW78zR++06ddyEk4luqLop9e6potXkpCxts0d+GEZtJTn2eMY
3M82PwfNBHXho9u/Iovz4uWMphe7PybV3wJ/kcb/kHtAy6Wy1egKYzbwfb5wRZb/Myu6UbjYJeNn
QjfHCjaxHfrSzpMeHFCOLUlN9tG/usM7zuC4u3xm0MsENT8NEvf+sYM+P4xWurUJkg0dnpBx0N1w
LvtT9oUTvH6gmPrWY+Ocykhr2/t3687x5SM84aoJE/g11RmwKBxmLOc969HZUohmN/Jw0o/79FDm
NJCDhRD/EJqbDJCspbTQ2I6Hcj7SdhwmZa0G79xxZkwdVBC2ZWc+AKm6hKtEKOGIg+Qf0RrdvDLD
BdOYW92rljC6KUOOQxesQsOhxqN6pgjVeKYGDN2iT47hEaGGm362U6kvRAKXKTFrfnjlX4hwXNY/
l3p0fp//m4JtgCjpzTMFolaybKLalwub+PC8oN6R4M2sjqrwXc/QVnqdK0rt0Xc4wH18+1M2g+0g
FiI95dh80FyyoirZ8gWVpmOa0vgVqteJ+3wG5YY1fUtDSpPhwf73WLUsN45D/zoiOdirRp5KJqwQ
lFDrOYH1B/kXmRDwGq8mpIYXBFgM7BVnLBu7CCTX2Rsem48SlhWgD3xXIshSQAl/7v0FLJDPxknH
ccoRrAmbCT+O75ACLm7KwkmSWDogAVL91++3h9AxlThs2eTEWHvf9tgXR7e9qtU14eCCPt2rcN4P
l2aLxmBWv+1yMs85LYRMtGraeztYoKM0IkSEC0Q9DVO4RGA80I12lu2UN5Ybqv/uLU+2b6tQDf0N
OIC3xTYXEf5G6JiSiLg04oKgzGn6/sYH73neNNr8Z2y+6e1ikl9oJ04HgQibqDOmoU8FNysvR9xA
Fc5uCcE5ZF/Q33DNdEUYETOHj98ZY88S2l6sALNyNFWM5XxD4NgPwITVGdHS7IYQkXg/Cy+N3nOP
UrHot7Gf6Z+CEWkwUo7MzE2n/sWL6No4Dt7IaHZ1sPPkYsHbO9z9R8QMHVfEp1/qUdcEeKCID26O
U23lUgck0HvkILshxND6OciZDlKlPptQyXyeJrm+pVJ0JS+mUU4J7fWvGILf9LLhXLO/JLkBRrOK
nqpl7lOvh/9JQTTznYxWod0Arc+z9sSgxL3NsTWrb/yVnFYPe6jzFhs3DYLupUhek1s04Rw7zi1A
Ci1w1fsxxnqUg8y7D9ds/1C/NTsEP0Jel2cC/bMCQuUIJGhmmXxwqUWvwhzXx5iS9FRqQL7m/Hy1
9OhGQnJ02fNNa9lXZQZVzB8gWr8AaatsLjTmlDvCdTmz5K0ptNDFwEUcihSdGZzTfSmR+uxEoZbF
GZ6pMdJvtrzt6JaVuhzIX0jhx6puO4Rm9FQGJIbVDfuAJiNrbAkhSNd5wR3UlzT5ysOCVXhnFHDt
bhZXkeVsKZxBlOTU08yimOwE/VHS3fbAm9S/LvYBZjjO4mE8ZUenCByLe0aq8Q2zxNJ/e4AnFpyc
e4QJstdvOO5rsdxdGWjbTg8VR3S20w1KXZKWDSs/XEmzi7EOom1L0D9y3Ccsmz+J6OW46KJrfuH8
dKluzJtiTrZXEj3s+Ql+E6vi/Ulsr/Y+by0ku3Ztk+0KkMi1V8v/ON2wvBPw507JdFyLIQFXqH3b
DrImxm/2bPLoc5Q1wX3+bYx1MzhfHthmLUSeVStzaSTrZosoedrgUNPIBZgyK/Vs8C9cRQEIJW7J
oKAZT+zOumLVKVIwPE6A1XoZUpr1S1q7WhpkBgkKHfqohs0e/C5s9Ldgx4BcKzTBUmhUVjuOaO/i
zHyJ6Lhwvxp8hAnymUb2R843dpxUgKlGboe+IHu+yYJNHDkrFd3tNd8npX0e0iL6TFAxq6OccFtz
YJ7VmstWguGTKmoBIcLHclFKBnPeu6sOf1MEsi5E7b7T8xxUBUH4kmtsK77z6zs62kL8niiyFFbr
oloW21R1QeUoLalwH2jl/4HRKS19N/ykpY1/NCMi1+OVG37VYtNLX25Zb3TS9Tr/BwIvuF60wBui
FKhymELKPxeZtsInu0dycvID15UyIH3bVeJn6w4B+ox69e0pS1EBwwv0LgRqeiM788+N9ofbUPwd
RWLG4q8Pao/0Id+J+LTL1Bep0p6PXb52egd87TpvPNwAbKvuivmeTEFGkLeq8eVgFi7U7h+tUhHt
HiThpzH/XVEPToo2gsgAx2ky+y9CtydRopt1tWnJBmBsLje7PhEmZsBgnZDjFmTGJW3iXKc+4g/e
nBAVdrNwN+GzyH/C9KKN0jja5j7XKb8WjIvSu53KnLLG/4jsnR3oM8N+ZuXlUhMQ1l8LBUZ2JIin
OMedCAigbR5iTPFk9y49UU9YO/HYodznNlGfhHCtLlFSnJPCxuUgQC5/qCj4M02BoP78yqO9JVoM
4Qtiuun305j1hm/4FjGsfDWoCcv45PrKcYjQe5hTKgXMpyIljJpBZOnHKmGWFxXyfxOKmt9gwYkP
7QJZI/uCTGIREWLrBUUdHDq+MzvKqLWlwV1pWiTFXMhgbP65ahGGpD7Fddm/Qqq9boM+9l9HfI/t
bsY9BqIsHM98cMct+EQWm9YfYZJvgT2WmU2KzshmgNL93SlcOcuRjEgCECW1Ce2QE9tWvvOnBsqv
D5MQSvo+zuHK7FLo+0btjfeToG9VgHHCh6j2oNB1DJe8bRu12Rt03cJ42Vxow6XrEqzQl5jA8Yhx
qwZIZYwfnzqgLbfoJSLRqeo09nK6sL1gfZ9myrpryBN2O3i88zhUOSkbPW4YjszQ8xBJpl5qGWuN
PLtFwdcanE6AZ3XOk2JRs76rBO1p+iupRYG8r/adHwNdTrUAqKgp/8vKbILkMsa6Mdnn82TDwN9j
PrKvY1WZnUaZtJSzGTMNZ35zQiIj2X/1fZCLu6CTp7YgVZz49s2C8zAekHWMWoSVictAoY57RIY5
V5KTh68OmeydOtvHD4dI2f9PRNi/6O+jyEiz8mBC6MImWAgi9p5TARXEX6SwHyr+MlTfjqDuAxxn
BeVAxgTuca9nGjQT1BYDsWer0T1aaaMEvyivGF4nkhgFBmNzBTcSfBLgCyxNnAqKcbC8L7HK4H2e
YzMeksH+CrCQYxOgEfC0wkdbecSGU6HoZ7NjiTY0LudAfIAIVwf1KjkzJx521vXxRwfORYDhaZQH
CP9a+6q1U4YvERTdvF4GGLr0vbyYEowwN5RBmxMAnTVv+zAVUU/d5YJJddyMtYEWB8+6vxaTwYLg
KMC4Er/lVeLhoDr9oPIFM2n6wxnwmekljwBhuETut00z+PPA49nORK+MSNgtx05w1sa7a92XTxwk
ejJD4pIpN4ZJjXlJGlaY8nW8ZOEp9/CX6QD+QKLFZV5XUZ75Nb8bmoi2FOAPjlL6MsBLzrLUbZ5S
gdQ1tgqntxsJ3DjCzWaPXHVLpvVRgITdJvarDk9joaoDsjG0EjWZjtJjtyk52qLxUsDlVeYSXXxA
2jUpF5tW4npeWcu10pdFxmSLMqNgVzuQqYm049CNemKz8thOgaDJVWRyOOjyf23vabvs0DgD7gsT
3J82g/Bt3T5e8OEyXbl2V3jxU/Eo/aCNRqtzxvlir4OQngvcVaKMixp1W+KdzTFvA6PRGgtldHi5
dzK4MeJP1IYJaLLINhuvmYXkGbXLdviDvEzdfZiY4j3hfvCsgD641lQzUAuFOx90dbHsmZtFbIZw
ab6Sj9b/biwb6PikDJmPDzlGETdGVZA+kXjyyURiSi3u39Lb9DVROUaeaAsHCseE/44DmKHZK31Z
txjKD3uKbgaEhH4JIxxTYPit36ME7V4QXR5hJtKAInnkXxe9cv5OwpfkEU891WOsjUfImtoMJG4u
5GSo+HdiN0gJt0Z3M5QLlQLgLmXsoSkxOJ47ukrqDmzwi7V6Wpa317Va+aQ23tRyeiQff5cU10TD
1ON2FLjTN4xqBxRqHOxct7BdGJjCc3+BXs1FfIve06ZVeNk/r9MFL2COzv09gvTCbtgPnyQprut0
dbiwSG9A4FW6Z8myFbtB1jPke9yTsULE+7gJEVlNI4DqVy8LbvSKygqUbj/wEIZ2kAEZ3kEAxKmH
IIuF1Y2q7ugpXimYEFaI9W5+SD7wsCh07HWI5P0TKdEX94a+9yTewFvhXu4dz7oMMasOe0Zq3kVh
7/xZWNN0mUglEoFZtXJizYQLlq4kulFf2iPLWqevxsXvFjCvcGIZG5+AFEXM47HF+B+bLEhARq0y
tAw7ZgWjjZVdHyNoOD+GiodpS327Ik1GX1WjZRMiFsDGWe3WFZdtutnqLYUAAWNvhkCNH3jYyVWi
ev9eVTaIX3D2vaIQ9nK/X/bg6TsYkS3OnT5+eI925ChIWtOUPD+gT6dXVWJjkzDcY6QngZtK/5Ab
ha+nO5RgHCGd48pbm98BRixzPilPnmS/S0Vk1zue7R4FoPt+qwXTjin6nAIVDgBe2L03FYGfRhHu
sPzVed5t6J6LFY+khLONRl5G4GbtS61frP6rSpSukxCgYA1MCtdSZofXRyxfo/BqMPevYF1/q4fd
qzlhA+NbjF1u2QeoHtS38TJyfUlBOxqEWpetn21S5aM5JVqQMiBkf3K+eiUoc9EWkpB26iE8kyvj
4uksvK1yHTNpthVte2RCLoQv4RPIQDvmPxP2JMHghFEQFFkXOiFkw6kutUHzuyowcrVoceENIe/f
VX+CrS4DUR44sePqIDD3FZruge/UBmEA6KRVWH0Y2CYbCqy29IIcS7kHt58RVThiBdRj7Bchcwmo
ROI1y9R0d8JT0eOHEvlx7MfyFeMCdNJDkSmkePDOEOJyvX7+UfMViGYfLohx9wciACLLpmUm/FB7
iI2jQLhei5Qbf7+0hbYKv8FN+j56O+GhfL47FsUc17qR4JcNk+P59MavOxRE0Sp3OhWGAuUFwP/L
TfGjlgvQY8LUCWmeZKyQVFKq2REja+bi73+1GoR2U00xlxRaziXWGdmWAK8mZZTEBE5u1OCSDs3D
BzSb6dA/QHuZnjYV+hLEhokXH3VO/BaHpqjZs8bVKxRChWgdiWH1ufy+zjrQ+q4ahNCGHv/ueiQA
TjkQIxfSo/CxWdK66EV/lpY54WT0bmOk8aKo/qv+BWDxEFqAZZyjFnbsmFxAJh0leetdRIksVgbQ
A2E9Ojpreg1KPYoZXvVCnfGhFN6uDqfNtU/IbQz0ytAk1oi7YUhLcXt6SIATfX7y4ZMBia/OLP2O
8muBnYWYpLr29wad3YKIIlvBeihhDPzNUoTrWahPbHNVMlFYti3q4jdqOPzbL0S8GxI+/w6/uHCW
SHaDu04OgiKRZ9PvJEBk4KW4bIiBcBpubFmDPpBrlxgHdLUaCVdXABZJK6SXZeQDKKnaVttLfTuK
jxYcSJC1RbcayCfU+I6NTHXCVE4K/ngCu/fnGXw8oMlJb1SWhFiB8hJ5fy4mvxPNePGyp/kszB+I
5R4AK/Rky53Pi1mUeU+mTgOqo0cbZH9c2AR60Pa9afqtlGkFgELLsw8qhnnNZdOzQ2opmbr4HHZM
UyueR4vZ6/ySx+JkvSK+Ox28GgN2afqWHU+HqfaCmvJ/9zuMnj9cAsir+8+6yR2i0BHkesYRNSdb
6wE1mqf/3EYyUiXB89y3koVXKkFWD+13Pbk3yO7OT88VxPT+rMf2NPfDHM5Id+P1dqnaYvEbkCHh
E3KT/ReRET0oKR55uuWgfaliMpP/asMQ9uFY3xHpKSitwmgyLGVOkUA4T8qE8SFNzpkg9wQ1YO0e
Pi98yGgs43HORwCfeqo8BjK3rcKgh19SesMnD7P7mUJphu+BUni5xTxl/8eJC1Rko85a8GU3vCe/
bZliEp5+5nmV9ThlK3816Wdz/xCRbBkgoLNp4FXu6pbg5q1ddCg3iGQnuYRyml9e5AcoN7F9WOrZ
je08LAnoi3U/vgZdm0T+HWE3l3GXUrg5aBkBA8f5fydg/Lzuh9j8tT56B/Gu1hvm1GSrfEVRxevb
+EBoTbIRYWzjPIhY6bA3j+YhC2XY5Pp1sD0+vNqrUXIE6/oNej6umhk4b16sWj3MzHTRqTj/g+5Q
b0QaT93cdfbaiTGfnUGSX+/naIYrFKNRR9eQg6vuXAJufvpTz2YsI3dK7rd5mauE2kfj2gKlfNWM
6gRYTr3J4FW6GhaA2aQr1Opnh7XoLbUaMoruJGtFNqh5cJabhWLrz1hOorVsbqIKvI4jSDtgbpyG
Px+xsnFlze/vMQrcnOgVcIpTZmn5hQ5pegjNn1bJKfL+pPn49uJvH93rOQFkU0KCTEX2+N1dZfsx
C/J0GQgoCg53poLErPBwNp+5sDsZGV9K6dpwGYukhxgLyIolbg8mkORwyHYXD/+buc4YTmXCDgYU
cqes0HfrJZ+XCcgupCexVhqGPL0PQrgyPVV/28+6ua4TYLaH/O+ESsirpaQcPCbMMktLiF2FbqdW
Qe13JmK0eD9KZ4yMqw2FOODkNDX+c0f6e5OjnhhkZk4WnyuUM01/4fO9IRndzwgWdy5RyUVpSCXc
0Au688Lhgw6qE4rt/eGEfCyIMaxptVta8YLmbeDF0WfDxsSAQqlgZFaga6rxPes5Y76FMIggvfsX
nZHPaMs+r7eRHn6R6s4vPO/SdUiecz86UHIFN/im4MejcvaHKZ8cdr1Hjs4mnGd+qlrINP6MBtkn
a/qmJVBzj3HNnuiFxjDCNXNLi/0/CIjialp5zLKeYroDZOA7L4cTAdIOwkssRbhslBpE4WYy/y6Z
Y2SVQj2B9w07qYlTvciKZcnKRXwwrtnaQkmIr+JaBQTDmRHgw7UjxYlTVedeljVwprvuj6vU9Cnh
43VctKLTm9HH0AHR2eu6hOBfyQX1TxQiIfk19/jYx0zHSsGK7aKToL9sqgnPKk9EUX0suCSHVx7Z
q1RiIuNdEj1Ec748kHWeBtYzIdkuPibkHdTaumQBoddVGoiVTQoDrD4c1sfA2l1pee6VKnri7aHl
ljlKwx6UzTX+ZVDyLyf/vGk9Lrqoil/NnaHwdfn4T7XZWmm/hrGhnaaiNkyKr0U5S9g0X2hPhSIQ
8xoSDyuoJi+ELq67neHjdqfFnVYb4yM5Zna+vc2o0He5GwTdITl9nwnawsfX/IFeagH3wxKj2gZy
I7vve6GPZ/kPvyoEl6whWSAyNetVrjTroksNICyhj6gvEBUP+eQPfDfua0ymnw6yP1gjKAep/4ru
xJsT7wGMmvyJVrCggL3QOQOzHv8b3jgwtZuxYUFXZPN1RpUC4Yi9eZGU4FAxjVvv+j1hWh3i2QcI
9Hg/75j9dtC81ZN77euuoe4k+au87tIW2YbS0isrDwvhMQDIoScSnSHCcyw4LL0N6JkNH6/AGjxf
Zkix5Jn3IudFDiS1Ah55O4FKKIHF7u4M8/aM+qalIzIjCujN6sGc9YuSMk02T/TOyKFJFD4r8s9m
7MglRsIQJTHppLFPM14T0bnFwujvt0kiFvvAJWE+O0TIRmMxYK8VodwmAHWIFK9n064ebIAu7auL
qxux90rMzgtr8pi8n4+WkDppyX2h94c//CI263vebn5pFxysvhzupGyFhuxo2IbG5a0vvRNbeQdS
jUDnZzCtLYlUljmfB1oGK0WWRAIi93Eu32VByB3U5oy4MhRQ34Pr5/6H00YNp1mxutkzbXCu0Utp
RHfIBN/kmm79+tL17PYjOs8EVYSINZep68nGyfvIYoP6CYWkkKqmcv5g7ZKco+ICwT6yj40TjzHU
8OURT3d/pfrH/3cEH2rj+hgyz4MVdKlr+Xo0BFTO3+QzVHKrEd3m+HDL1rH6mKQARcU0w8Jjzasz
PJvLgv6NxHxkxkVBluVF9hLHnDH0PtOtqQzH838J+yQkpZj6UI+CxpVawTc5caxp7A/wCqbmj2sP
2VNt7JSL5ez6HxZGH/+yq2pU0wRFWpC1Cm2hTpApKf1h/gl6m5iBsJSV7QMQhhM3HQLdzLkp7JJs
xthU6BI+5kwre69/6UDsSafizEP9sjaLazlOfH6BCxRQ0V9OjmLiWSYO6XCVIYE6gE2LBvQdrU3p
Ga/UJmPtCEf4lSe/+MLMTMwz5oCm2OnIrDWrHBa7FKFF4QG/H9FOW23x94wV1n1dQ0l++ZqPzig9
rPQ6EZmH7NlgzKlYnjzSjo/8T/sOWpxrKWcNQiWVuvldZBSr+efm7g9SOhfXIFt9ptVpwwDbUCgD
AZ7P0MwD220FLQK4mVUzfuKtGGx4ROTavScR62aSz4yd5SwmQj+NsA8fNr0mIJSFUlf/gtMGNrCY
5Skjo23HQRzYgujKtZndygYzvpBUJkKp6YG/2c8OWYJxAxkXidRGRmT7/qzw8BVAr9jHwEyyHFIs
zaCrKZfMReWGGUBBds3iGV7H66VDXdM9b2ZodD7th9Ib/EcgqU/AJFepxzzSpGokaMPB0jXDwoAv
cdd+pEWTnc6YggHT/fxje1clldO9LpQV3RjHQwRqn7THRQ/GG/D3YU2bg7rWTO5IuGkRFo/zud4C
KAx2KvQBFzOG+wOaBI1aHd9ILg6rGKSE9JleZ6J5GBvbij8+w4ugtqGV+J5mcnUovwzzwgd1XROj
OrzkggQNrml2nvhjD2NEcShH/QkM6IAf972WzjyxgtI6ojyWQkkll+Xei2Npggq2Ef479nE+GBNE
LKTBwc1W2olxb4+jBk4BlfgbQjOq3gaWxJcvNTZgFHY5hmmVVUXAuJSyDvpoDLmCSZydpiO09aZn
Hrb9qp+vkbXc7tzBHJa/pGwR+bg7lmlehPVPsAtB2jT9NsmcYpZ9Ifw6Ty/Ybahl25XLfGIWSjrS
9FcsoOovvl9yiIAB9VPvaETC19Mq9pNJuhlhqCclmMLyw4aBvRwdT2hISgVB8qtIDgWgEopLVbri
c9nS6p0qqAmoBQkfx2ahROSR+3fOY8SlFf9FS8up5x2By4UlL0+t3Ys35YBu6uXL7X8xjYeyrLNY
jH5Vn34qJ7d9Nk0N1PLnH1cfUuPsw6KchI4jsvdEiPDXGqwxvPHuEADFIyAAA8n67bbZismZ1YTJ
8uC+kEclHTQsyn1jNXwMWuibJ8zux4u62bPv3rl+IxjoYA2b4kOYULcddECSrQ1otfzW1ml4euNn
k5EsWJAh6xhMwEAyIFNN3VbmlSJTOv8J2rYwosi22JNGJgAJhYf3X9qlMCtMKp3H9/laltIPw5gc
mXrNhiZMFt1aJLN/H49aqT8bpkuQJdvaCFY5ZTR9W1Kgct5y5nH0qqTQL8qfPLoqKi+Kx6AnNZHu
rRb9bgs1ZqHyKrd1eqWyuPm0bMCk3LKfkWVNHC0Yh3A/QdZIt01kOgoxT2br1fwSPQDdcwJDcsCC
ydjTyJGAEH+SWky4j7GQtPPwrFIBoa/ICzeyaPE1W9JO9ZiAuihFpHguBS1NRc9F0OpjUzxBNj6C
M3iRRtH/ZW2bS6HVc1FtDD8U4dLZAHqKpUGthxxREOtG7rlSNyAQGlkZBirLZoRX5+FUfs++/QaF
5/lznCIKumX2IX2CkFh+NLkk15MZzcwKgezGqpwlPqYEGQbXEKH1Md366434gqXK5TDNlMMyMWoz
Yw9hk+3Ry29oUGX7N/TSy0qhJ1I7Nn9ZlmF2gm8lGf1WAMSLyt6MjyR1tf+q3sDI9fOB6nAexZ7I
J+plj+GQhGraMWXSJahiKG7bpwh/gngyuf2s/HF/6vZSNmqXnWvIZBWtVd345Tj/2vMpPFBm5Xcv
u61XCt8lTVbyUz3yZQDesAo+NUbAbhhB1BN/9a4S0ih+dTM+VLtDBSk7v+fLNS10DCF+qNQVyzab
aZtWYOM3gAGlZR/JW8smHlPZa1YcQyCcc2ZraKHCRb04BtbJRP1o1DwO89j2YDI+3x2jWyfFX4SK
EzKZ+2JKPpT0+ZmfBvtSaHuKj8cNTc+ZWxIWML4wm2wzisifGUgZIWiidR8QJMl2HQCLbtZUcFse
wUyx0ZOha1z8+K3oPRQiBfhiTTW4fLQu7Mn2HiJ2Ib/wTyJz9rnnkhH0xat9sx6Gi6VcXuu7SMDa
EeMd2BB/w+SZ9JRtyKPDeVHbbBYAQaNDpB+v/VFPrHkRguiAQGjOgFe9QQ4A1iRY/6nOKMs4HEgI
C710cpuJ6fkG6bgv0j5DPWL4DjVpqpzPagyDDogW2tp9aCEQneTH4V5y5RQShVpR783CqSrJfqGI
quLx+TePva3+OBJ5NLnJ4XHAREiHHjY47ew/0TntD2q/h8wyoG4W8366tw6TM6so1wtVZy4BgVq+
bMj5g5IZN9xqNUsuCZXYsfqsO2/eBrobt84pqqfqLZN7lIyltRjnH13J18zMLGp1pU4zHWTRrI7U
I0V9WyizGdnHWP0SwP/23huy65wGIeMy7yH4eP1jFZJy84LvZqfC/0dAjB0IGGetU3UcD5pPxoWG
PbRLd4nt+gsMsWkQBgFUlS8DVeQA5i2PW/2+Pqv6WYO6PwBPG+jNKjL3EQgvCgX0iLUpx86tpCBS
uox+wkHF2tUKtWK28AA2p+ozprIFw1sxk4Wv1yGxjO6r5dIzFxMbBWRBACUkMZr4xuAVTNS5AMOq
iOr4Nr65O9fP8EikYtqMPnv1YMxECz1lHCyjgsD69LRYOabgHLtVbO2uKiOmttz3gOYwhMO5Cebo
RTZq1CrzOdJa15hxM0gX77ise1qc52fXv71VEX3pKSOjBTkEFXNKDeBxxCXkyX5BIHRA6ySOGBHU
cjF8KbEa9fPWjXkOMo3tMigCPfYxdney9bZIfqnfqXRTOlo9Eevn3y3aDjPwEQEiUxHwvOOe6yea
LIEbjKC9ERCUzEPY9aMjIVUJEvYn0Bcm0Si3iV3ouGKX1rWZ+Y7LJouRuE0XP8bjh6DwOiW+swQ1
o7esau32xIFhAo+WtIv8ysfxG05bkAvKWeFsNSxj8EoNBpdQvz1w/Wg8tCcvDAghPfg7oFiUdpvG
fMbIi8zLx6S98cUrbPKxG+ISSNdytl0HRNAfw+ZksyrkaeN9cCIpZkqTei3xdCXSZ8ObFWb1uHgw
63UqBveO0/XUXAk5gsUCr730oJ2kCwhzoYmIKFykew+upKTytOwH9hMeS8pOtQU527rqIM+fF6ef
XHpmwwzgj1CTdQVxf2eMcNGJGmgmPyLsEBCLsMVk/VBQoczsqT2nRg06CXNBBo0bW+2URXoY0Zci
TN8xjCGG1QXO7njDlFHN2CrJUkipDRUIWS7giWIGkQub9pofEBrKX31pUOfDmKsV7rkQPfY9FoOJ
rSnXNyq7xrrTCsbupoFaapkeMxgD3/TmV3mQQO0RG1ieLAGgK9oGv3X05jjNeKLt1SfSIc/5tE/Y
QwVUrOqW8Ox/jYO/lt6ckFRLLx0JRr6ykXyD3zwCkbWRO/uuUE1TWOZmDmj1Hl/cBfTlEvXqKWX4
Cdg0+hjiKvBo/zditk+mYmCDWF7VyalwbV2etHBqe47IHVeX5m0Wwkf52TdlD45I09svUJelAnm2
dhBZlMziZTxze5yUp9EjYFU5eu8h/62aTPtVKN+AkS7+nX910H8HKiL5SkgbLjSAeHuzowiSQOeQ
VIvPRTL8o6Ds7ZXzSwbIDcsVT47qT6iHfxMhxd6cawL0o7kgpMmuKiGUOE0Ys/UIxxoLE1VOoPBA
I5xrYu65kYN5z/Gk5LE94szIhW/6EB/kxdZAefV/xAMRRYZbF+jLhw796Lvx5rjpdHGWqIkiAsIh
3moBR6wKPy73Tq0huG/pIyg2tyxWL+Cvs9NmEAIkl4JuGiEc+Ju6H7NeikFglngD8pSMkxwD7XBy
LNoXO5ol7/zdjI0WtDMZRdqiJ2J1/U8qtdHYmRnzBC0yTnsY4UAlzs/1+Pw5xZiE/IzeHva8/dNX
MgWtQJEhQ3xCjJGvRNUoITzC7OPjHxozGav8AZCWy2/WtLWWwcQMN4gaLgEn56fmbDCfxyi1Swnc
TnWDmzb/Q2dc7lMpTwWmc5jHv52bhj/N9XKyujL6vsaDslmqEvRzNe2iourhAE9kxw2kN2NBNarm
xt4X/57VNxU6ljuQg2ncplDu44ANh8ig47Ji50CgxtoNhIMTdzMDswa993ql4lYWo03sLjXAYtG3
uwQqG8uRZxE2CxKzzX5rsaANC80T13UL7x/T1YzDMSxkb5f849kGJh+pGfHZTrNlQAyWI/MFv5QT
cITtnjCTtcYY955IGq2BJSo0RbjETRlfcJJH+WAZxErzYmktiWbRTaOltQ8XAZYl5jHtjb2kle4M
lDkI9NXlbRoGl6+LRLsvfWLCHYMw/CAcUoRQFw78ZSy99oibKa8AlC4u6sDcbK02SjloePoC2Q+E
XcU5+EuyxQXAC9YWk7BENYTukMGZ1SerT12OmwUx9qA77SH7eXZflskMOypFmBNBQ+LGqxyy1IHi
RqBvlsBJ5c1OcG3+hoy5zmHpQAGB0y8b0bUG3Mo7BqsRfUFxYRMXqa87A3YumoUVuKhPDyO+yDHc
arG4SPiTWT6rv9/bi4LcJBfKLdX8MFoWL4JBqSqPadNHfoq04wO5PNfDUbTX5mjfRkoTFSMb5xdT
wHgqgfpU2DsaXAzDGWqvpWtaS1pFVF7VlqPHR7bpYqVAJueD51CHugXtP9ISNrZ7pKUA5VCT7TH3
l6xLMOEEi13VBUACFHvYt9sELg9TyD3/rUiH/c5Aqqt3LxhWnf+a7utdXPuILDMvA2Ah/khzcEWK
0z4MKQCxztCQrhELdTt8JhD/bcaCa8EFC13TWH9ZV9rfkVGo/2rPyZ/HT4IH+PNMea5GW7oIJCv8
F/NHXZH3SK7o0BV75+q4swguUZ1NU9gt1JUHozD/W/TeFkijqvEQ9mVoT1qmgyeVr4DqTL7YBeAB
VICp5WxZ4jeVZP4z1CYTMccwGxpGd+Qe0w/WF+RQonExObswc8bnYy6WOmk1llniTHF+gF65utUN
cpGWXsB38rb10LA5hb6h9HeAIXMLW/9slvFZgefMW+AygHEu0MYZfjzQdGSd1Tgb5rad1KQSLymx
Yp+LyN1AqvuRjcc8B/+uyad3iIe6GPxBYEeSWyH+MuEtdEkqINjeD36ojBbodoVEgTDQVy4VFI35
pscy37c2vyN+zaukuVifuj/4Nu5IIamrcdROtGkTxdEBL4UoafQcPNzxUzycnMQLcSe1TkXjLtzr
YonDNv5p/txI1JWd/O70+ugr6SV475TmFpdtGbH/lWMuWBGgxiYweyz0bt6XWaoohCWAps4QkV4h
LQzmvKUNAbEpJ2LND0AH9rBYaNBuYZJIDnxRrlhVmH6dkqplKxEqBBxgGxHXnJxS08Zy8xwkys7f
Q8/wCPAs3Nyh+nh3kh/NwvItKLrA2fiiMz0HzTuAw/3UBC419jvW+2TthVNsHkdTJOFT62RqE+yU
uppIiGxdLigfF+QGdJsdp3aBYq5ri1TRk9uqKtdoiT2WYD0ehCWxmUJh8l+A17k/AYifDVvyAh4c
fH1+AyHKLaD7n1UzZ+M6fwbYoBjldX4sqZUGOUfIVyCR57cy55z2E2dg9EnydCzojHLfij/Le9hk
y86sDC8GYm4SovxHOQMa2J2JAf+iziGtoKUnmUhpyH/HNd3ZDVLvGOdekCrN0+bBS3dW+uHekFtQ
RajJsf7kwoFENHR0sNQl4LS6o+gD5rJdE4bZ5YyOO9xK4p1qpjl1Z2u6Hvb5yzoT04NVRHUKXLj9
YDJL3FHCQKc5ET8OzWeIXXeO0PlULKpaAMa7qfEvwSpzXeNFDkJ9hX2WhB5FeXBXVZv0YJq57WKc
1+Y7YXAccuqeIlhjJ2u7ByRi0uMTDK2iBpbk846BznoX3vpk/A2NoMG5xNv/rn7HVArkDfwC0x5D
D3pbXmFmkL5E7xHh25f5k4UCViw2ICCdtfJ5/dK7Xpl0oSBRPcn/w9lUgti5xVzFgEF1CjZrEzR0
o4YyX7YEhTjFIGFspuJHdK6nmXLyNAHAqIZUoRf184Oo9DZVunw0pyrKIlbW8rJKVSJlx4fSrCCr
okYfesxgeUwBJrSLIbZD0RIit2kzaNd7rky8yPge9M7Bml7XaJjXLKEz3RhFhMIGQa4UdIiGOM0P
QyC+N2dUU4VZF7dYZcY38FWvrPyW4xqxjyF+jc1XPCCUJEG44PJEz5VGxhlCcl9YOiiGT52+G4xS
C/nTM6aTlwMDAEwD8yvp+w8e1j6GOBzDDm0C3H0ggkcs5SfY2UJ8C3TN4aXReT3tT828cg3h/d6L
6XJOHf0GeT4BfsjiyKr5wwOPbbD0yUobLpzM8lC5y4vpO3ovM/gJbRHzjh//iLbdL03tVWodvpho
9PSXitwNedOodVGib1zuXa1M7VbkYEhkt54xmfOHUwqUg04lkqn322EUlM+Uqgh2HqfNyGXa/qSW
zyDpFE5ZEp4W2wfel4iH6uZEf1EqNO6TvggA4N0mPOBIWgllFz74kKXxzzXboX7Hwynu6vh7llTS
PmWYeZrmvpHrUVSH3+NABMNPaG8PUYnSKsADNa5dHaxkot6vUUyVj058qA/ZtOLIde5chT+/sxgn
MRSx8QQ48UHDKQ44Y9DgOcbuF+mwS3truIML3egN8ImAuHQLgISXyBCf5OLmgEjixhVVUAS0CH+Q
AEwDdrlWv/BYKTXCl9BNS4pxP317vmqxvpgaHd4NJu6MC+IeZ6yyHPeqWjdA9Ioldz0MY3mxW+dA
Nd35KpiRTT86C2mEW0fS1DBJ11gFSxGt6Fy/AmJ9tKK5mbdqVAo26y2Vh1SQ94de0r0A+/pnN8Ei
md1EOJ8SwMOIdxY+TYRHCaQExc8Et7ZKT9a5yXZoAo58QhDWu8t0y3KNB20u4jTN19Yv3SgR8eXj
jVRjN6a/yVwY+y0uMqq75vKwOd9UOb4mZEcNt9M89oyvj8IxQtXJ97dzdozRpSRl6uPm47asgtvE
d5IBDye1OPr4jiQLt4/J+gisHLdUbY0wN8c/ULO+Nz3OIXITtey4mzclry5CMC18wviZoqE+MKZh
2qJs7QH5pOe49Bn2pntMasTBIcfLu3qcbcpnK33qe8Ki/Sk772OB7tD1rmESLM0PJPrcAzI7WTI9
V4Dly1EuWiZSdcqIZiu2/W2aP/09KVCfNXD7fnGuUilrT9c2J3bPqTBpmyEbgS87bQAA9bPTnjYz
96Gd8t5WHU0F+x8kTMHd77eIXx/FvGnF/pFTpXAWjoBef1GIcJmWI6DOGPM+AZbEjiXLldURp6IK
q8ZZkJaH1RbqAWIpVYpyyNLfC7u4g5skVLihI2SClcGR/WE2uoo4jfRpanS5Bi0mxuhfL/fx0aZH
o/lnT1RE7m+kmiyCzjcAelbSiI97DN3kZoCRB1vP8cGMPsKyNXMAxBHYgiVmKewtYjPtG51Abuwr
jajAtYtrVn0fsCkTjSRrNINBxstSFr48XSDTUdrlqRwWsBkJJqwvrYpRbHAIw5Dj8/t5ArNrHjHc
V9PGtQfzeOQwZeTBuWA1ycw9rTe36H7YNPdsopWFaY9z/xTpBwA2pPM8rdLq4nOIUKMKgVfXMfvy
eMn/+8z2FQqNEOMEivmQsChxn6gi+KhxwyoeeVMvVQsZ6LrotfxPn9T715K18VUrrcGd9sxnEdFY
AsgVe3DpcAFg5nq5Zv0FcRJ/0h35Ff0moY0OuQ2+bKPtwwf4knewadi6BxGAbSokYU9x1s2pWa4x
rcdWNngiBKWcXlzkoM0jcjTl/EHL1CK0MHR1OL79aPdNerqoNWL9CJKEzg0IYxBr1pdqP/UmqEyY
TsybpVbj1CfML2zXNyX5Xzgbs1/zs/k4g05vsWoUdFY6RokueXsTOOY5YXep+BIWSLgW1FPoHMku
iMO5TZfJQixgoLphH++hYKfutJNz7GwvoC02KtSiEptr66uTRaRFumxyYUjz2GlrKONtjsGQ4xqd
deJjm1vTbOZMHfhJ0aKYTVGC1HMldfdRcqCfcDoEq1Er5m1OXhuWlUmeirru9rE8Pw07jiXkMlcD
ezO2zi4zs1/1jPqedjqnBJ+wC0zJY+lF36Fukpy1X9VbbCOR5sPoUyuCZW+35ICw7NBJgYyDrL/n
t4uKLIWM9NnYOHGHapkR9lbJWH225Bf1bh/ceLPJc6TKhR6k/Zj3qUTgOaeNYzWsDJ9w9wTfdMs4
eMCH227m6x8E8jLW+P5nFxtTUsnHo342q3/rROoroDcwfgxAGLP2kQ+9rDUsRtv9RVUAUcFNCjNm
BDPsZD0T+g0yMjTWo7PuqX1cJJO/SJgtZGYw2OCrW5VEWMKSdHaWBP8FstPx5nPo74M6WcznRVV6
noK8WyADsY/y9fHto1ngnLkKHbTxW69FJZJYXit1V6U64ApJV/lf/juUqHC90CtyUuuJiftqTHZ1
22/6Pwjo1GgeSSIxSavxeulBNdS0q/1u3Adx3svC/9K2AJEgTHF3z8K5ZsKUeJuJqgwJqHQBScBT
7Da8w8GGiBbWId2m1pGGem0E9xFoKbTejMu1e3WS2+5W6wZmnqP5EaRF6ZODuc1hlZwTF7cmj2sL
iGc3Sf7zvA0AJF1f2SYwYqQEXlTSYA9ngn8xaeIKCOipcshrPDxZYXlBfDSIiYAQQCMGmY9zo9aS
F3AI9bng/n0c5waP3eeFyic0ZUlAUth1/U84/CtyU8fPZU92/XUvub+TpDBI/koOvZN2RzUV1NjS
KnrXO83ebK5Fvi4d3odTTIMWhrlLn922Zjn5bN99ZzVtLGIIGUu8fltJjRucPmD9+G7iYAnzDvC2
Xj6vhIkT9SDiO1fslAC3SIc3ctdpPE0POu5+g9p63zddRIxgUN3FjJMSqYL+gOVhE5UuC1ST1zxk
CGOtTRvNuWkmD3dcfBWx06nayBzZTWNQAWJ25lEKAlMLSX2gySBHfiQgZbRhvfS4mVA2V/POuKqI
+f0h+JMUy3hsbQbbHJS42F8MxlWSTVgWtZR6gg0LVpDg0PpRbMSbbZInCDgeFhquGTJagBmbdFee
Tz/PahdHJ3nMRfgXlhCk8Fno5A13ceq8OavpAQV8yg833OCEH0gA832jSdUxTPTmMqqPaImzU72R
WcGjQVSN6zg785XC3M46gbeymn/AGBkizMqtllroIyGZT6XKR02Bp3j0GNOVLeeytR5lYH9mghpD
XDP/S7cV/zHyaH6QG4tP+WasBBwc+2Qdeu8aycDKHjoxEd6k+ejb/WMKo24CvZz48LSm0qzhMvRX
60PPIxU740QBYgdGVe/r9AVDDdNSfholkRADxHKWa2QnlOgDyeyFmGsPc7+1vgmWEqg1qA9xjvDd
lgsc7HJzvI+2tEXYR4Dr37btEAZR60ZLhpA3V4q8RNuTtju3tTEUfURhA6xeLMA+YoJC7fH2w4HM
vRgZrnP6y3CeSWcXv+WUGpQcz/b/2XU7B1HVjDvXx2GBtxfPuJMs2XsIgouT6gkaiHYa85CM6V5Q
NQmPmibDb/khHPQdBDnsDLBS5ToGHihsA7CCJdTUT1lV7nODubjjEKiyVFfQsNcAiDO4WjERxc7W
VzISM+ekj5YFdfeQkZg2cDxvAW0uBVXi05hNTLmwOMpmFJCY1Rb4QUAvGVPcXD/vwLlfMN8rrspA
mHP/qVRJ57V62M8rjorgcIkuujVkuBoPbsWOmdB9mKSbQT9t3C0Fkag0N8W/WXlZsUhslPxXJtNK
47lX/QTwy16ImftsPBXLO897sb2DHH/y440JzilPb6F0hyXOWdx1bQrG2VecZ4lIi3vBK1vCw0mR
k0HHxdNu2h3qMSocKTfylgGNOr3YcCumZsGs2h7JB3E8li1/MfRmrayOWK8v9oI5kl7XVaaaxyjU
Vlbz/0pYoCez5FU/CQF11uzTM1uLCF6s1zKhzOCkFSMCNzEFzMzDTq4ULWqLlR1s0AMSHeysuUkr
0vzadLJS6oSCFvS1jzr3wFm/9RKHSEVDzJbzmWAU8+cTYzcGvOqqvOf+8UmUpvUMfdanAuPnxW4d
VvCl18MQfPKueRLSabg1DcC6LJ/qV1xR7VKNG64c+9WBrmmHElwCAM+I7Nkbg53Flc4S9111QltO
aEnQOJ/+Nl8AIlDUJeht4TlQHgHsTHlzqEXt/VHNt7dz6vaoz1dB26lJkjoer/OEs4rz1oi6q9pn
Guc073hp8wzWmKg84w1OwzV24gyQyLtlO9y7la791ct/qhF2DaPAzSPw2Fw406iOdbfz2ncWmw2/
fn5KLZ5eUEFZE/ounRpm1bey5xhTA+7J0yyYxqpQisDkCm+DXUkOFIB+CoX+p/H9jh44fJyh+pGU
FCsu6skJdAy2U/ZCWs73QfODQzucQK0G8kZm1bD6xkBS+lD5g75OdAUOuQ7CQKVqlIdSo4l9tOlu
RsaMIef2EEKj4zMTDv0fHgmEFYz7fqTVUu+VyyXs2INf0EkgdYi0PlA4IwGW81kGfeAAlXGJE/x7
mFvj3O1JuBby3THzJRM+iX1DcpBalw7Sg+RaY+0j0y3v9EqP9DGbgmvoBkhQbbrD6bbtTdMyywbI
f187NAkj49h4P5TU1NokLTF2UUF9kiDRHwUxIRQUNGbkhw+Da0Tt5n3YzpUVT9A6VKmyGYN2h0Sd
ntG6wJouJ0nYXUdVBh9BFgzrfdR49LAJnnfjL9OO55iRMv72A9KxrswDApjrhhBDpK0dQW8dqD6g
N1fSBzmljM2NPVU1wpJ7CgB1tpJbBDZ7eIQfXvx9+7axTbP0G2qiT7fqxkYNpEplUHf9JV/0BY6h
AkVMD8lb59VqYY6YPFp6HIX8ZjFBNUoVxuor5wW+cr4iwsZfYfiN6ZtrtiUDyq/Z/mKTFaNbbBST
3Z01EckKKdBf+B/LYeYNJdrcEujhlu5J1+kj7JpJLToYRk1RFxXySVB5RLVO3ap+KEnY90bGnixd
QxwNLo0UodWvrEbxuDX0H4W+9ojZzc5FZzSKVHzcw/yjQx1E44/OySTLt+7QUAHVUgs+k1ecrmgF
9POvJqeIE+NCf/hYRsZvjtbG3Lx4tTgSnroeuQ+DQhsirQRCkaNXuXViaEZV/k+CMfqVRZyTLFeA
ONyCgWpDv1jbPh3URkbQVIr0RmdpGgyp0UelRpRXLgKu2azB/I3fkmOEyzqTU2xxwwo8SIGjfFM0
Lyn9uX3sBVBXCfRlFGsoeq7C3Kta8DkjEvM0QdgfuVULBr9yi3OoqnWEzrpgtgNV13yKlOnmBqzk
8pihoIGfB81iLMe35SWk50YZVtCYoZJ38jz91+R0INFCYwf+AQO4PDBSpaj/2mGWpM0R6VgVO34o
WT9APRfs3q1+lT2x1t+oNaUTHNxAUKxweLiEA8Dm6rAZasXM+7Pd78xyFgDiYu/sLLG9T7mfHsHR
BA6MfADa/H+g7vgzSd509FWUcpG4mPs6xdEjGLk3k//nMRrpdokNc+JWsr9PNgWChhOvjQqaupWN
/T0eTTVFnKbjizEtlQxrPG5Itn54hZTlGqsdlepFlUPlcNCgyDaWv8pdav1SlvP95swneAlgbLVn
7M9qcLfG6487cEqdd1PrVKWlO2En/KjZVE2xwpyb86880aHrq4NLrZeEhiII2EwF4jm4qshorwKE
9kbPXDeagQXA4wPCFos+JUTCXQ1HSdkUmhggAwfKIVhqAm6lLjI9fcVtKutYLuV5YW5ujYMEeU06
9t0RRzcKAXQTAbw4Lf9T8PicEaF9Tvd2VMF7txA+cy6cfC++1Znd0f4Mpq1SwiDS6Ztr4KWxuBOp
PSMqgq/RFp6NenqIMH9WHTiHQUpoUbmZXU1KZiR/JbI84UaJ5cgPjHpGgtBCgTntwh3vZFzV6BCj
RZRoI6+mzqOlO+3JISguU+Mf/ArTOJddDNOKYVNEN4sKT4juuTcM6Zxsbe2M9LpW+5CiPJnzKt8r
IpRjAvhW/PEEQ5sVOtlhuIncoNIV89l9KApLKw1DRprLx6/LkrDRgNfSnZ+LxAQUNC887HXcCzQZ
mxCNoy7PJV0n/VoIRA2U9mx2hmZptqdJMxe9ReEs7UztewjoUjLVbW+w4jXeI8LpE0lCJektAZ9e
Pg/IEJe7aprOBpWUQij+OOVa8+fjoszbF/cfMR7VRU+jywSDhahOX/LCohLPSlwlsa3QIeDgdCtj
Z3aKdAVqmLb/Kp4pIA8LBkW5UV0OW+qa17/wXfp75kruOOCPK3Tr5AHP7prhEU961YNQrW/e1+NV
zVfmK/QqcEtNr+7JOz+3jpHNc+/pXWKMfI6L2DoWuawfyKKXyUA0cuTXRDHVFTB+z05mLV5kyJ1e
MSZynpqYp29hQdIumyjfPRHZ8NuIMERkwY4htpuPGWOxcbOfTVz30wQSInNAu5UmUb3sjuZUTgFj
i0tuWFykpNLe3xgSImykKIGAzNbBV9nLvhTK9TTGPR66CCFuJPgkYdcsZb8VdjL60h4Zm2GG53v5
UyJvMeSn3svBqraR1SnusSXDtmahtqL4gQF0Wex354CRncLcI+dijJ5L65jHOuJLL+hPiVExU+NI
XvTGmIP5kkzX6E7w+P+EAua+KXCcj5Y+RMuFKCr1rhhYEKAAoYc/gkjFUkbdvOvs/AnIAME3Cyj1
NUMt+UE5odoOMo/j8a2X/s00netIgqX/OO2O8LiSSxkstg+GLLqmKOFwgcmlOkzmA5+kqL9CTUA2
OJAKalciX/rzqzHKbULSWtsV890GOP92g8070+2gr7T7gnWqmFyh8zBfYFqoz7gO3hum8xjooQrU
zZaXl+wwQyuwA8owghieyKShHYUUmez7yjwXhkg4/oBinOPX9y8Avj4Nnb3HAjT8pCC1ruEA2sqE
YzRo9/w0ED7erjTAeuUIymW0O/7KOG8IDEWaThF/MsxnHcXysUIK2IrWOWH+S0tsZVDPMMAR/TGZ
Jf/dxOFrC493LIAKNAOF5ji8qbDzCWP3zIItPxO63cEDqTp5tJfE4emlp543mkwIGtJAuwIusvU5
CrbczUiF35bw+J1dxr/3ZBa2KyiTs5T0thuDpxCpzyt/BmwST3+OsilVPWga0eZswXssWBTY7S+4
f9TjNHvBOSSGE6BaQXuG0jg45wYwAFPLhKq/cruvwHnlTJ2RJmOF7mRU6KdXoCq3bsvXGIVRz6UR
MXbL7Ge33nnS1XLOkuWYPzUzysSnFp1YEU9pykF4gzrnb1x4Qm91598tbc03IM5l4GTYXDAtQ9hU
70q540YwP0qHDdo0ZlwBRqF5UvJj5M9r9oMLJgftvvfZFw2mcBLYoQLdir2CrebwI7/buZjMJPYW
V6oIq+OoKtg/lORrBmDMoJb6a5H0vjihBlf2bVVcGgwhVgZlLx86BiOPJG1UvVGE5n9OtwoAxVx9
pZ1aFr8gHV488uWxANtXNE1f8zWnyHb2YsqYIqocBKnXz0W2BxBN1ZDpFVwWVXB8RtHV65bzEucb
b6IS+j/gP1attYSf1V03pvU/wRKYW1WTEosS5OPfg1OX6p6l22dHf3mGvucoUzJp9KhTFmECFhpA
AmuNSqc7FIZjmSzWdDMt83r6kWy3A3qLUgdyBoap7haOhLff5uHrkgbdQTIUE//TTIbpomj2ESbh
Gwk0Iu8JOnWUNoo+GzAeL4eFY6fWhuZbxEzREZfujXFcV0DlV0P4TzNOAtIdATq2R6rAN/U+4z19
bSf+zh04IiUjZtq3MMnMCuaSRLmXn15PJvCRSQryhQSH4j0tkQn2gX2guX/ueb1R4z9ic8jfB48j
WkbPPi9gDlKInDS9mAIAYelpc8+LDqfoACWvtCzwVTgc9jL3105OtvG1F09m9rDZJRpOZ57q6ZKt
0nCmtDOpw+LRbY6tUelfzBu2/TGd5fndKilPNVIrXOFhuFuavoNyHiMeDft3L4JxxgNlvW4aBcOZ
odM014Y4LzdszzU3uNFLrXll9Eh77EaNtkOGDb8nas+rKJF7cySenVDxbYh0WkIDuO03tgxpX+Xi
t9dhiDTy0tjqPyOX4ukdxePBqMfrzVih9aXVn/RHft47TPvcls9P5o+t4aSvljv9RmyZkA65qACp
LXeLA7bEfXbCC/v75jnqflKAHcG/QVVcosS7Aopp+8IgJ75dmoUt8Dlqp5flEe5RmpCUZ/fQE83Q
jcZDRym7mh9/vemBT6wvlT1lU66JE9PLJsm5BMrNtIAU9Ioe+joWOg0Bxy3CF2nMxvDps68moxxj
EqP5uQ+f16hoGMc5cqZRsELlX3QKTKPRBv0aqqrHxZMyNrzQVrhLAhp60qE7pmojoaAe4+ktnZtk
9jVoQYFpRdqKMbjMFa1aGE0XYDjAFS3kT/1qVJdTc/wxt90TtYus4wp27KHZFTdRU1sKFmXDruZ6
aFSd1AciwhTN3nIm+LYpuDBX32td5911utRgMCASPoeIz4yupg/FTeQdT8hrJN8scr/4u082B+6r
jhOct78aB/XV7IB0levEuBYt4jibMpDq8kv151M3W+wl7BK95mBWSJ5HKhDEwCdDk+V7yygt4yeH
rqsHKA3D7/ldzDYndHMeatniZuVELPl9RUKJZoJDMMdSZGEEoj6cmeGiScSUbnUOH15hIzR3qWh0
Cybzxe3ipm7xUP4NyST7Wtmd/YznPzCLqgSmoCS7CEDLR8qsQPn645RoNYd7XtSsstA/Oj6Obhoe
fKQlM2A6VSepBbZx1rabidBdSsrWk8o0Xse9gZ+V22UlrDb9vA2W87BVqtTexljC5R0MAHxRIbDA
FLy7gR8htd1c3zwbHEt+Hb5zAHFYZ8AZAP4n1Zu7VgowLDD/HwqOelsKt12FOkW5Jxg+/cdFaexy
9f8labGhpgsy9lzKbnf45tIQaShXmmzKfY8QybbL86FIUBpoAYfPaiaQojQH5y98ERX2QYT77UjA
S5kzM6ZhA7dwAigSaNL0Kmn9QfVgkqO5w9ZN5K8lKLZ4bEBTuXqdPnTDT8/ByFqaw7tPTrozofZa
7maRWuYhAm5LA+tpowvFJ6hUW3VOI9SIqWA5shdeQv2YU01F/QeKljnBxWLktpxZdjdznBrKqRFt
8UvUXAAbOy+GDHeNjNdCMdhBjBYVRWe4kaBUqFKs5tc9wfetrZM/T4SB3PobH6vuzqT9hshzaekj
50nh1miYhJvXAOZo6JnGSIvIXlRNxH1JJYuALEqko0CGqTNGe+K8RKatQMSS2twckKywofxnE4Qh
4TVfaL0SkKVlL7mK5HUWAcQfBP2v1qP9yFWwpvGC3VXIq/TA2gWwjHwZReI94akkfNlyEL5rlvzT
k3chr42eJ6+AB6kjVppc6wxN5lj6fvxkCaQxVD4pg1tYX1LZ8RztmxQJHKRjTs0QIXYTLe8XYPth
YxK4ewOGmeF+KLE0iCtOaK7a1qdNNKHjUP4gQq/lNyhKFnx1ybx2gdlmVrlOjm1sWpfM9Hh35hvK
p7SB8SFt11Nimhxah/jUcs5bacRfRN7iRFtw6stWmaUo4/VunxT/O6Dq0Uy8pceBGgU8IH6g5GxU
Pq3EwurmMp3RZN1xvTDq8uFXF4M0fvxR/bWbnbuXHWKSMgM03PxkSrgPg3HfMcqX61IeHEwYRxpV
zbYXqZp70iN94676mErMr4h+zGfCTbKro3tFS37uxZRgI/AhfAqhl1y5055GO4w1Yz1GqMGpV5l2
tMtOtzHW2sAmJyyLasZ3DM64c+t7xiXQdMzJrVs22ajFiIyYMEAZycXaL8OVdF53PyS5zLmtzG8i
ArayL+UA27c+dBN3goMYxGZkahBK3hDMo+on26KUYsWkO1cVwrs86a4ERx7rRTCGrEG+4t5TJ4b3
9Az2Qdxsjrqn+T9TozER0307yCer1RVKmYELenuRWQnJMqflRuhkzUc+3oXuNImbFhgJ3j2HWf3a
3ws97O1lL2haqWAEAmLJq1f/Q7T+ToKEw6/fonCs5LBWo4BNFdj66ZLnlynAoJKPzPTIGHuZdVBC
I5laqq6jbj4OAoLEAbzkZN1SAfW8ZSuaXd7zjG08dGKA1t5i9xLxEQvUIJmP154ZdLNuGWUbKT+Y
QizfGT9J/hC0UiQIxKNZ/9d75739kOS2DfP2TtwEBg6MXUC3Rl5SYa7RrfxtejGdQM5C2x3xs9D8
fc2apTtSTSCMsV9YkyuL31JJCmn/92W4a5YHjcbW4mFH8jWd6dyj+01H60aYmxFgXy2ofiqkAmnf
IWwLkkV+pIQshtQmwoHJSrOpG7UGVXFD/Zj0eW5WkseTV9+GzHxZUhr/mKVVYaEQ4mWQ0SaGOzjv
13cF2kOsG1+O8hyqNy3ax6Pc+LhsbedJPhGxoEccxMDBe1qXyNHcyDMfjyvD2/tVwobbMyCKIlX4
pVvuvHnYxNnK5uCEqhPcUQJc+yDQn4oZmrfRJb03bkPSFaOgKYOULDn+UOnoyYhI+M053QNVGeRB
PvX8PfKVMzLlrwg0aS/FTy92Cp20H9LScdkcyMnNrKdSKwvYNGl+GhOJlIqb5HZEF4jq+seU20Bw
tawcHG4176GX6NkmdvfDoDOyLApeOt1gnv9p6yb0D4JrZgoM4HsTmHMR9yRT7TTm8oBh9og6B6Zt
PuLD/A10XDqVyJJszSoIzsLBWKLGni/US7xsfRHw4o++sOQCArXAOnhypOTmRMfijIEsq1NA9Kin
sH2CctfBgs6XTtzigdyOBLxtFBtmcyu3g3QBva/dmJIux+Kx8leUG56I4iAWjenOSw2Nu+5bDw+n
hXg0WzWaWb767MUXGseoOMHrvOUaxOuJUTxATfMqtw9tpmd6rBXQafCGVm0SArO8ne4NBw9e6vlw
xzb8V9Aa/oscAZDeIpQiU0YFA4JsfDaxuNluZhvF1GvTUz6hkZzHDVq44kdo2t0qk6YGtrS9ZyHb
ZOQqYXA39AorfVFbqoyNE4wwTcJPTIs5p/FS7jxp7qZXFNIHm4mycI0OQm/rQjYBkjLKqX4Yio+2
uIS+drBIJQ7WUdH3M9pST+lqbQ2PpiMCBktNVYGyjDd4YhJPn3w91M0P17MbQgCHWLf79cPnSepG
REZnjjFosy/EWpi0dKJrXJAyyBjh/bIPBoK1Zh95q/f349LDTQj/o04KwMV6Ezb3IZ96c0EuYa7x
Lvd58wEydZyV5ZUSuRJTEQHJ5j70h3CCEdceV8FW1uEV+4h82PNEF+fYw9YIRk81QxbxRIRLLshW
+a8LFVQW4bC6/0bQzPcqpZ73w9ilNQobJ2iUlhCiQvET2tnbA5+plTfrWy+qeBYWU0EAzYX9OujN
B2V3xNWCQDHvTQx6XFDXvczXsuC2WTdt4JaeU9z7lBR4KuwkTIVr8hLaKbuJ7Yw3UgcRZ2jyK5W/
OPcw4kpqr2RSLKMcKwwNecPrUaomRpGxdPrBN9eZxKIrh8wihr8sUid4ZoTWf7728Fg325L0hK6a
LSADb53rpvTXfn+cifu7nLizfsuMkxs37l5XQIaermu32TEs8okYrN46R36seCDGTalm6MAJCJVB
RR0F1VfdnsL0Yw7AfqSeYQgFSrwnSMqrEEphbOgY4m4oLISU2lDDIAiInTFvGvcjP/a3+K0FMhnz
SOS+OvDFVLLWkruX5rrYEG804j5BfInfCwU9W5RqD1SEbp1K4NYHaVPbAQkU3wjxnIiORzSgiB78
ND/mzlyRDNTprs80FpNLx9A5pZqusSSwV2tgA9OS7JDLMl7jrPooOhPSPAtbMt+TkGsUdiMitqlW
vpDMTYZRpiUGva84SDtz/PJCFIc0N8tBstsq8tpm1HymKlI3wwfB6HHHh2yOkU+y/DULP/8CjBao
2ZTY0mjgfUw8/Wp75rTUD70p1i17DM9h6nelXrqe7wuuKCuWg9/L4hGPDFKznVwAsyB8cnaIV/Tp
j6/XilorqbwZNcHLyPet+2XReObB8XG1A6SKaRCQ12lBFa/JhvqQLpoxYgQ/qnUwK9YIRiCbmYoU
5cJnghDxWw8orLs1bqT7QLFSaTlIFnD3ITTdJhASZaUn+08/aA+2MK9X8swGDBaub/2TK5ICxOSl
IWHmezasmYsakP1O9sXAWiiFryos0krFCYIlYhI/SW3SlQiv0Jt8DTZLWxmjvLdHFxEQUnS2oze2
7zWM9g15G4tMOuoz8eyhbIB979Bi3VONmBLVtUEKcXSRyRQbmSscPZj+R7EVimQcQut9wg6OLULI
nVRbbgRYcsD6/EgEKV6TakEumXl17VSjHnF4H0R5QGCsa+qF481i0tIHr1t3IyPqJKOPdR0tgeQ0
zHlVVKoP5uS5Jqs/v9UtqOej7/P7JtVTH+fQYcUBzyyvMvzebZpvYxRtQQBoefQ+XUWsZMlIkOtX
qnzMT8YIXyQ47RcZbG8AwzAUrCDgDCOGVP0NTHOB6fhpO9HNTCYj+YflAq09YRW+K030P2d3zA9V
N9cDOLabgkMJxwdtZhygvIZUf06VyH5tEFcKcUW+EptPKkYzIdFxOecTU6VxTt4EA+Neh9151w3z
s29610apV9vrVCOkYcysIJwOM9c+MQleobsdyIRrILxCfnvbce3DWAt6sSlP9//Vuh8rz+5SNAkB
kTrB/AC7U3zapLA8i5ccEYdBxxHDc+JVMmtQY6y0Z55z9aFLPKPDo5NHNyMViUriDwXdPBrkE9sV
kq+IAWgGhJWCOSrOo0Wmw4PuchqfFkahRdoD35ifqaueZS/3skiRkKoH7EuVtjEDkbJZDOFbODnG
UZNQ2Iiv9hCW02LX/EJEDasQpIY4m4FWdzxGUSgVex/8lzJSEnDxJKlva8b5e+zo0/qWfQr0Rzpg
ah0RX1it3weUItKXsHPcYy/Yy7+0rpqoR8uxF5GifjHJPJT8CFafxgKYy0HWjSjehBp8dWuxmwoR
K5lHo/D5LbYil+31CNl7GHXJdKT1B3K0b3pE3VgY5iIIo7nKbBPVAN5z4d7dEaCTlOk4Gf7jwfeQ
WLtD17K8LWWDTqXx5Aml+27uJ9V7yFQl467jNxkPdqjN4OhonFP/lZqkxSD/PD97oRsD5uSTR/VG
nBwVw3teVGy4NiqdEMjcj4WvB3hKmzXFxtGlTUvVU/+2iSIINIApOw1pbPJs1EQr+5Wh9B/CkkTI
ANSYUuyBS94kQYDjACx55p/rnigGMgGuaY3aLVvL5tq+TSowKj5t1R9S2LRsv1nZmj4bilJHp4wo
X86JcuOBfAbLlihRmYQe+v2VqSRAAdnGQwQn4EXwfqutyBfXlKUca8dF9DaNMYdJHHcKK/hWVF8n
NvhMbfCF8rcHrwcCLcJW5HcylOFQwGcga6+RsTWfsal4Xwa0K8c9bGCPFZg45AW7H2+PyjR1uDRa
1r0bualyQ3UfZUCvverthZcNGoKOeVtZKms8qAf1KKUQQxp8COXKQvq4tc4vojUtTWGft0s8Wpxa
thwwzmKGfLARAYZk9kkuGsr7cvAH6L89IiCG8qmUnXroQR8AlNfJK8sKZJmPdNqkpM5hm3vD7KRg
E5tZGsxP/lkULYUigGwhaeiwF+32tNKG+LEUeT88l7TB25ZNruqzIBnmlppILVYhGCgWQmcfcnsH
8qgy8EYbLiT+6yDUovO02jN4Lf0WP5fepQ/kDyeL9x8NFVI2/1zebDxzDKBWxzwe6I/tYx2753VC
kxCxn6Gbcg0QNRLueta8JgMvx9x0A3Kh85910dJMqFY9GzkPMPf3bzOKPba11Nhc+g3xvKeWdghx
6+5Y20oSFgahDcNxjSnP/cKzHGHDuw+FHIC3eb8FYDL+62ExPTTu+U9QIpikSrWlQvv+FnKrs5Pp
pIsB0nJMeuS+bSLiRmKas0ISjSW4WDvnLy8Qd2W0u0nEhEZmyK23k0wCqdOvOaUZTB5aCCwROU6i
w/fIJsQEN2yTa62IJnMv27kmmpF3g5wdaynjvspJK3MR/zmxM1WU6Xvkhlsq4Hj8tbUunLXVcL+z
/kBUxL9qXwoj5uvrrmZo0SkLYSXqyPIPTYwTKl/2YSy8nDD2O7BPbmUQjv5kC/dvJyrAXKRHeLfb
9ysPEIsrfzqzmtXyOfJZbZZKNDyuAcJ8iPwz/Pem9GOZ0Sc4pQmUQHzwYGBsgDc0sen6bkgCot8E
hPWu2cXBlo1mao27sRCmALHPwVHu/sCYlO/qh4n5epVM0zPEwoOqy2+34frg1lqJSeATtjSNcJFE
fpsqtkyvOCBlPqANuDf8P59bz/aV+xLpMy+COoOKnOQGrZSk9dSADxgdkLMAGzj/fk6LWv9DlF9S
4iOb0bYAAulOgWao70iy5e8/WIZ2xaViitVfpFZ9bA49vfKoU1MM3YHCHvJfqfPm2/5ycm7WEveZ
cUaV4BfzbCKbOedU1VRi6KpW/tIXFJXU2nc4514RNao73/T4Fdqz8YG6cLtkaEHCznc0PvibFnZl
MSKq6P030jeJC4ODGEL/189c2fUWTOyEwU0n3ym8GBjrPPBHR40fMf4mVDHl5hsFCNRUXjCMRAmo
TsgkJP7o68KPTEv+hsKlrWf4IRRgXHEmxYRMqRtd346PhoL7QF5QQTqo3be8CvRdJpxd9Imfv044
JXQdjAMrCYiX6w/U1HO1ypztQaHVgPx7zcVzvWMlt+XkstfcYAKIfM6AzSMWa4sfuEoVxMgPrLDI
v+/L2/+q9VYlFIn9j36IAEWbIexjj2gAMG2wFiuqBHvuXyUzyPG2HfEZwho9NqyTm2lEECiVY6TI
rP5voM4Be8uxyIo4Yg8d/YUF7jen44ay2jt8dG6xE1GsTcx7PmctrsFZ+leBn33XD1Du8pGzefNV
z7MaFyI9gS1PaggkyCO07VgK8Re7Fp3cmw2jb16+kgpuGVvkKzo0duleGHHrshttahIv1HFfO9LM
Zfhn6ZGnN++EhP+VLdW8a8Q0wRuE6BZPfZnC3weR/blPsbM/yMklQebWmCkip7prVMAX/ucjsYfM
gCgefiSP4ry8YXpG+qUSu9RQfZKTGKuo23Oc6HHKQGKhwxi7Rs5zkjKrt6eJtFybLW8KFfyd8G0Z
0URWg8pCdgRnLQ49VxoT0aWsZat4NaFb+vxBTy9fzMEGkib4/6mrhZrEUCD47kt2C4FBGTlR8pkk
jx0F3N8uumJNPqrHlBJh55u+j0NZrGTYIVMc/sb2hDGKYJ6MOajtoUBojE5sVbzsjcgZ0JMejNKK
CkEQNsJrjjh44NKsVl2qcjfhAaHDeEWeYc9eMyLrmTSAXXILxTRYuL+zA8kAWtRn0+K/dMH2PmKJ
Uyr0kjihN60RHaXQVCWqquUXwwc+eGqEy7PZkIdCuUBx0XzDoTkJZjLACOl9zCw8rui2zc1yqkzm
DKJ/4NdsHRYo+TXMTHe+RnUMyXOCmfDcY2GZhP9gsXIn0o54Mz33oBmlXw35PkUEmqrM9zXswUpS
Qv4IC23LQCQe9mMRWRnIIp8YmaxlZUXwqNAJY9Im7vyB4BApIjhGkdep0wXUCzqw3rKpO00c5cch
yQm57ZQfP8mXyr6e4fz/kqhsb5UTgTyFcmhEiG6XhGkXzBcPbFGy010idGzMBxtPgk8imY2PWcHe
xAVudmtOhFuftnvPBQGLWt5PFt206iOJ1zkEk4EAyj6yw0h6lKHIobxcDehZDAAIRGUKntn/JhCc
OJv2wAMHe+W1NEl3Et+3AHYDlyInWuWWhh5Uplv0lBNGb2rbIqD18sYCOtIdTI4TSmgpblg//GGU
K/zeyOqbTM50JRl+4TDOy39DFA+zjR1+LDIjiImq2hifX6e8Hu/A/RvszjnftpwmMRd3dzINhQUm
0EfhorkybzkTK6X+m1qqq75V1TMSGdKS9080A27WaxyOfMqskaLKTouKfj/M+W1JLi9Xr2mtkxtb
0ZqqgViHX3gEKh5zQuHfDS0c0tGPnOYavLI1inX7Op25+acj8v1jTBP642kMkTUBPGZX+14ve6gi
e37bUTMHtLZq6p6k7Y2+u6Kj5quTTx3it3bYUr7MkjGUTuQ6CbxIyMBn31bGG/JDExPiYXbDpvTB
MIjT16nuOogC2zsIlNXyGQE315jS18t3B7RyXVKAuqm9kcRqWQGG/KAeGNvv7CEDUbBhKRWA3KNT
5iUYcwzep3opz+LziHf0tm2RBv0nP1EEwmzC8o6li0HuMQseJbH5s4hAK5qbmjWaG+3KtUhoLx9d
ufi1qVYJtqrpGed9H3dpGuJn8zDtHeMW1o8hSgEX65klHXCDg7jkkRme7xSiPOlG7ncTgbREo7EM
cRDBO7/89Uchsv6ZCaJoiktOKDQ32QHaZe1WIRS4eqAfb/0wTC2F46QzClF9y3SLbaBj/ZXzrwzV
HFKQQu+JtP/xi6VdNpAXHRxI8Lj5n00022s7unTroiuvDxK1BUeNYd0Tw7tmtJE4jGN5dv8jMNAC
EN1vOib459vkOzid/8kdx9+cuV0ccw5UM7WKMulJ8Pa4KrBVZQojkZKJIzODn7pLwaKesEtwMiaa
IzZ3jr4+0x0aHJ/xKIgSs56ayp2tM4pZjAwgGu8Crm27Qr9DPibXjnnGuELPU49Pmqx2vXKregop
BkoUTTQHLfg74B1W/Cpp6CBC/NHHzpzd+Z8KsLF8NwjfjgoZYcS77u3ZZi0Q9p5ZCsQVQrG2IWrY
GW+3kOOqNszzgJRaoyQVzr3uHDB+fZnuIgH7v12iJTpPyOmBgOp6PrULLmcHhtAJMvvWQM9K1NcE
ztUfioUYVHzfPEJsHB4lmJ2v8a2J8rD37zixWqWQ+MTYHO5xGWgMWs5Qp0kvdAT5XTsRvVnn+sE/
dDRzzTbPR9UnYHMD13lAWtC2nOlSi3mJ8Ktz30PWNgIM8omTOzh/VBUiHeGWeLUKloWLor4IrASK
uZOmICO8kN3bwMjBRpgXN7V98C6xsAoYI/nXh989/kPwcxPYM46zQ7Xz9D27eYJoBzfnuMOyjPtB
g/KFXYSmcnTEdCPL7UnxxXqSAEg13TjV+yUwg78xa+ixr7UbnYsl7ruiq5ZdlmYN+psd2rhb+v1R
u5vGzUtxZcPkNCbIlRXnpAmFuyNLxPWehQiTPLIRSFO54ITZeUW2EyapL0+3YGeK5ChutSUyERWJ
oJkd+NR+ZWQOaUV5E68Wjr3vBJw5/u8T+f1G70/G8eiBAwd/IQrsmIRIZ2NFWBVFd2WTLrzWhZR8
0lzcC1ujqEV/tJyWbTe9Jspc5x2qwLkesLHRLK8ynofsvWZ5YRnXckd5fF87CdMRDCmJQUWFwp7S
PRQoO5mGDTRm7vodh9TIvCiCwWpcrBSHh4yfi5YvasqqD2ia2MFxwl9GQyK6dow4Nvav33NqyePR
2RPIVm3FIfRGsc3pI0WF/MARZRZThhmBPoCoakFwRujOdNSdIN3qTdZ5Ieimgk9iICFNa+cIo6wK
rRPP3Z+4CIUbuzFGMm6vCM9vCr9CratlHAIAc/U5B8uKwpNlnSS2nXJiK+2ggfL7cgGWHd8zCzAb
PTueN/NFtJ9PaRptSk4g8Su0rfhQdV4oLmkeIHjpvOwMrsrpczOoRfppLPEuLjfujSJrwsaZGHBG
rWrQ0zTdrsTqGp6pMQ9mVHc6kXqTd/mbRRYP3KnR2NNZFFbLVGYwDVH2NM3zvg5BbRtq6q90AzFc
2ihIHzG3of6uUcC1RXUwauYEbLyZzxp0CM6FRcsKtUiErGTQN46I+hoyi2tz8ctf1ihYBVTdRusg
+EpHzXZ42tpbb42qGtFTdCOHf8WJea0nmVbLlEvWrduiuD6qCAG5op2+WObjazp955k+enan7uzX
Oa8iI38RjGKojRxfx4Yowjku41DV+m+O7oUG9Vg8AFR/YXplt5zZijbT4VHxIzvpVBRjbEfAQS9z
SCtkqh7LisocBWQ4jtpE4wbNAcWkt1mUSYStiapjrpStZzfRY4PeVtOF1pYUY+4X0bQX1bBk750z
S1lwMFrT1WvmdYrcbZroq+bumsDIPpESFmlafLn6XS1ORFLMkMuUUp9jsKcPViDi3CSVv0Ne4yUk
g6JupLQ6lnRJnQXSep5N72sQey40qgihzOqUlVhTmY8WYi+v4v5X2nUYYM5NAqxK3hJWggAyfhAt
OkQl3w21ElzfXww21ggeXkHCiby5yGm/6jlfWCQyBnNlL0XXJOUpAcHCp1YXeXQ96pb33XyjBlgP
Pot1ftnSEKgzoeXc5E3IREy60Eb3Inr+jVWWIHpkmR13c9hyEsVWpcAJUfp1Gxv18mJp+JtJb313
I2NWKMeFbrGOQDAdVwE7sl/OZAtjVG4vMuTtOkiB5pUDHmdfCy1b04bC6xgqP/ZiIUQfEeW4jSOJ
4csaIlEXzZKT3Kn/gsV0XNua8d2P229RU/ka08x9TC5qmk3lIGxJZUEG7Pmsx3qJPOKv6886rPBy
2Ab08bISKQkWs6zKjsskXAjk48bwIvEeoMOhoTYjUmfAq9/5ZfoPFUekBsut7C2Va16V5fYiV2Du
KqpwQXjhGOgJYLiOMZ91JIvpz4rYXks609xMEpIz3+YB01RSWeVAchX4ltfX8SorwyS2ZeHBcLdR
oLzFYG7M+W/8TfpimmbDHZv2ZjP11XiY4wKYBeeKE/uiyy238W7/tjm498fYnZ3ZCaoZJIVqEuLX
sTSbkvWDQ9YW+W/2PWCJLpF9cNnWFrRDPPolrNPNOi0qEUjhkF+yR1Az+c+W08mibrginD0aZUYh
67q0zkiVAkMEIOy+B/h8pAnNMdICbFHlm/kck4cvbz6HMzn3i4DfM80/I03AiRhlP8uBsNxiWKhk
0P5p1zKLb0rxVPV5CPsLFMPdQykh1g+Xr63dk5PAZrdNyNt8uboBiGeoeD444wB3RPozUnIuFS4m
Ok6GtFM10lBp4mlkYfqkjj0eMLZrp+96jYKzZcazTXeVVlI69GTaJY639v+T6Mx3NQOAimE7+VuU
phiTchENDOEJZIbc0LzSDoZ1u9lfv69+/nCnP9fdXrwuy8Hb6Ou88iWc9/oqYaHkRuxNBTpRRBVd
PwFjMRFqdS+iT+wKnq54G4wq2HKGqecHtNQ+cxIj22vHr0WNdCr2kg1mrW/WflGsTtEakXS9xfTJ
WKqXGbcX6G+xgRjVPEdx9TNfEyQrPfBnMXmnMpYmOucu0Ys4byYw577V8MIdPdCTJgi6qHZUin/p
lNia5aVo/EJgfQeym3IgLuu0UHO/oYfJgnm3h8o+j50+s+IR9BWuqFedW90DFlIbmUlj2e2e5RMf
GvOu8SWYX0Txe9jMkftah/BcgeAqzdAY0YKNkzi5X9QUzhMawJ8ZCIBRiAqD9027RRFC1THx3lpR
VAkLshcjGMoBcsEZvPvgbZ43I59NcJYQjKNzddbo7vZXjDs6XyMW15HbgUxMmszX+c3idqjde0Az
flcg0IbDxQWezoaW9zoW7zyWlAi0TOcAg3Ol0+9EarCTX/Ap54priwzJyRun6SGbeJJvNvUCJNt7
kC3NGWnRCmTJBuX6bZs1WUQH52arImHefSA5WCfh3xc4Oe3Zz2M6nBhzZG4UoQjgBw8DvQ0I5qMv
W2iSt5wrkVh+PSOr7GUMyj/+ffoBT/YDEcyZMagTF00xXPWnDB9WcgwKFpF2g1cQfae+DM1jEsY4
4HsxW2EK2udBbVZCMfALUbYAROFov5m76aMX4TRN1B4YnNeXG8nx5S5S+76FGHvbWq9920pXlcqf
h4jmmgXLWKmhLK7UaHxhgqoOKJeCalInw/462KfGTCsyxc1OPOpZ51Rb/lldnFaSVqHw/JLz/ZCP
2VOr5mSYlnU24jLqe8mVB+r9eSsQrfr9e5qSCwGywAMkP6KTtQCFsw1olq40cRgv/Yu3rPnZbHBP
yek5qNghQebRcsPSD9XE4PNry6WtTjHEMIELwkWxjCNMkQE9dk4ka2ZSSDJzdtY6s4Mqe4QEB2Z+
fwFnE2u4wWfxOUD7Me4m5gEVV6PV9kERn84gRj0yVLBgp561hLbhBbUqbHXF2cpiXTGYXyhXo7vS
iM41X//nQ+huT2UbgMxohEa7Cmxd/NFXekxyMHxZvsv5F9temKsMarrQGr53vq1oZSQOfqMTSyM6
kB8Ae0nD3uT5efVXWd+7fvfKAeQ1OV4l5UHY5iChOd6lKS/995u9fBN3IGZJ7xgqAlVeRQ076UHZ
f5S4gXGkw+loXLG3diOtGtFwBG1pUD4PUVL99gB4ENxd8bFGrUU9P2TBQpTNwXQ5OSaXyx8kAkq3
IqN6eXMK3YOkiBqx//XB1R3gQwsPzBtLJykJoLKqEDNlWGfGWQ/XtXLwEUzhYq3sCva93/TUHHSm
Rwec23mRVvOwf8tZm6nrNqDzMd32TWy4J6Uyf2Z+z9+KWkQPO0gQiTdfLuZIYyhkR/C4Hc7NNelC
uXW+7QORD2yAK1nBdOWfwVi5MGEOAY9yUMXREchOi7fQ2ixJ9p+SZ8qmL5ZTBPUfKvgiYCkJaffH
AtcGYFhI+FB/ZUSKeCwNpMJx5mpC5wDP2VZ5JQjsGe8TTlUG8pI6S+cnZiWNPrpMrZDHEEkfQDga
iYnsOGooyPQPGPybFlzN5y8EWoXz1wPrQlmsZhv5qk7jqDi9fpd2FUf5zVcBYJ9F+h2HCdrhq/o9
WQpT+nyfPdj3gt9gtmhBjp9+Nge3HgQfIDCZAHLRAKvrwEX1Qj/ePYey4oVhihUkRbTli5MDg8pw
zNZlonhKDSFBJR4bhKESh8wPQFeWKekIdypY1qBldZJOUp9xgLf7tlUytuxwU2yvM0pdpghnWLae
39BYv0X3d1bAhCOzNr2kYBX1BMNIuOf1/LfAp6WyCetxb9Ytmbg07tqW4NcqTLJrWeLcmtJEsMU9
BJQeV1pLoeTDvB13lbb51KVjQKJeTfJwcnrMd8ZmNl80BQhuqYYEyH++c1rbA832liEyLZ4fYWZo
3AcUQmXqOhdPd0m3lgWriYZDoRaMhP5AtGd9xsokoHObMWgi0opgvgaEW4Uilc+Dggs03BsgDLXV
Bk1U9WxCISr+EQ5B5Oi5344XPC3mL8TLyK2QNR2g3t0HAeQWMjn6VasBNeVdBUR7QIOSsRk/ON2w
DKNDBn4bQF6JSw4IfAqQsCk4Xxx/hmrFTHxUgWDGNRL/sE1Y/8ErN7vyEcunD+S2U6BiGh46QziB
6HYVHfq2nw0eStK/bcvOVBg2W3Z6pOVDtcKh4pXpqbTbR9iOLCW3YaDCFs7UWuOAmlRdyn9Dtfi8
b+RhJK3gsYkEa/uIkeF6mpkUfBVEW2aTveRw9l59aFT7sgsuASLC3KPtrZP+fXTVfIc0hDgWv8Pd
RkJLztMfenFsNCqTxz2kCzetb3BShbBnFwzfQkaOjjzmEqS9SNcm/4RCQLrW+0WNEqQacnhMH8sL
dDeifARxXkiF2RarOGAxlncAWLyLkWCK3aJYDqJrA6vtc0i/VQJ3iERQDfvqOdm4hBpqQPf+eDsH
+zD0d1dSnxxhi8Xvqc0sho2J5S03NkaiOc+MxGJcDMmHnJxvQi7M12PCT3I9rAxKN2f7B+Llw3z3
oLAqXQM4t9zX3kzraVg2EKatNCFS5nRhU/NAMNHYzpQ+61qNPaYWkHu+XM66EugfxBL4iiFfMEmw
6SZGXhvE2oyMFbVddx4Qdcm5IMdkOQjb/ETXJYR4sHduMPctg2XZrdK/NTJnsG2xlGL0tyFF0z8+
zuF/3qXwQpHLQBQzv6FoTMKTdFM3kufl+9iue3oGkZz4IZU7cXnm4afQCOud5CwP15hacORP9fKV
RB+Z2WhxkRUi0V+dt+GIEy92647YXtSuJmBEppALTJHQ3vocA9kuiOASLgpKBtGexs7/xWpcUTHg
CZcbYfdkk3X5Xbz8EgcvP/wsU0TB23iWCy2Ay5QXbZK5P1lvXLUcvPmV+FegwcryYLslQZUn6eJd
JJoCGLsBoq/Keo5jxUkvCwoSueXEEmG3zP/lzONRP5AzJVf5+UlalIgqF+wg2MtTVmbTDPpvoRvi
JyRESaYksLoyDypSpOA2yvaw4bJB5CS3QFx+z/V5Bq3BbhlbvmPqOZ1RSvMFZToGT2k2erYIHEB2
Ttay2wetHMv18NWpHyHgp6l2x6+uRWBCt/t0X6tXXRBuMKLRZYhQDbC66pxYn6KbLIN1zof61foS
GjC2luXGalQswjEno/2IPZE1DHzZY1sXrmJLxf5/NDjIjMGO8tXx4PB1cdXYzdTx3fre32PDr1Ry
WTOAvPw+t7U13vM81oeftuglZ1O4rNvKoYpszU/oXn5E73yyzClLH+NvtT9spyH7L6ItB286Pekz
rZH92jRvm68WbzHUOWNCQ69Ym86YEOalf5yiRDTAT3FB/8C7sUSkdfg/AEwsRRqVRvw07pqTFjGx
8QEm/TuoNviTLuVCKMNCFejncTgMUGsFYrez9EU/gVZzNoLlQswniCJARMyRxknK/Z0SCfvtgZVT
FB9F5YTUrVQlVeqe+7P66QyG6T+JWJOh41wM7sxomvgbBlQG+9lviVOV5tE0LOsauw6d/bkzk/2g
Jik0xg7dromo3bIsAO1ozd4z2ugqBuYPcGy8zLTwjW775nY0JCGAawvzLwxvy6tI88nFUdjxDS4h
PYnm9zlQ1QI6JcXdDZnPV25Z8ofjpGmihV5KM07rWCwsaUO/OZdaJYbZUvuk8I64oMwnpP4nsrwy
kE+sD2Hdd4+WyaWIvxyI976mjY5DCpKLwibLZM9RY2WB6EZt3mAKVOj+/sM0z61ztyBmv4qT8OyM
kXgHD+Eq5vLEB8ZMhCXRo/bBXq1ypDMvf/S/z5GzTH9ei4/K8+XNJxqOUZGonx9pQ9Vt3C+zKFeO
omX7gJfnljF6eTXEsuRj0hnB7gz5YPRPcr6DH2Hyt13xJKsBhY0/xECmzbVlcca8OzSCcMmR//Tz
22xuIdrFfFqQaRf21Ra8bsiW4olyZGLTOHFLgOCsbGZJ5rogiij31rjpNhihWPTXbMgHelgXLeeQ
SoLgwMK/2ZB3uw9PoTlv3Rz4/iPrWmeL4ApyKGSGlsYJTEe0RecNzaBYBFdCyEBQA3GbkvahXp1W
osgNxvNX7DOu4Aq8Vv423t62g1b5nFpz7lwNV5A991mnUjzM8du0HnB8JEP1gb2yo+Vi5wkVC1y8
aSPXzxg5qkdE+1tzVv1t+YvZXIsU88z/wRaq1AIvqlXOvgKsUfV9wYzc4UKrKXjBloazjldrhdtA
4dPmo8EPp6Ik3BN3QQMnKR7FxiotRnF0yKPoGMJPyNidMYok6pKdXw19WWDadTC/UjHORRW8vgGe
fx+q89ao6pOHXDR4SMdr4OPk7AudPngAYundfR4X2OJd+FnvsCAhOyUf3hoJl3CPm9IngX610hS4
k5edhUCTzakhUbiZ+/9HcGniN7NG0eFXbty4hLFqIt1zMYAhkhO05ufFQRu9DpFVj9WlsbuFAwTo
d7LQdRSTSSbPG4A9uko3PR11674oa+jE8jhjp8ZjNK6a1YU3keGE4NvRQF3TiQ/oJIrfA28SMGr8
Pklgb35uVy6P4FmFaQ94BuuQJDVqBCi1vi+HeM4d53FFDtPcAHViSLxP5TE159aIJldt/RLQj/xe
Lfsyo5KJrzv26xgw5UW5dv/cee9lN4/DaEDMaChbaL73Lf5I7rLr6z5SvV9jAcMd6mKdDm4ZdAH6
X7skCVv/cnyV7Lk5sYqfqyKeisL/fw98V0VxSWWq33NmjKRAYmqmVKq3IknndyyIr2fxE1b1Mc/3
4ZbmbT33RfErzVVY3GiziUnAhsPOo7nJEc+irdUJ/sSlJtGX1T/wcAqejTR7MZDU7ZQ7n+gQKxSw
JW7YwJ/fCvw6bUVQwoEpDxnn6Y4dv0TNfj6JXsa4HyW7YDrhgzJvAt9WTVXvAfg/d+Ru4xZBoGir
HrCIgyy++esXGJjC2QNLDHSfHybeoiAdUQYn5IyN2NO2uLrCVqfGEbKVccRcv4pkYkyjF4TxJZzF
EA+lvrZjIXHvAbUuZkp4N/WYFns6/of3jQ3ScXPjQTTWvNL3aczDZmOhJN/fUrZ2zWX+zcpUYKPB
wb0GE29RmDZv2h6sgt2T4JPosaE+wOGTRp132S5D7fEoYgxJF5MhRG94EA79QxlqEl/3Ol4vpLRN
ke49HgTEXdgfddyF/WzAXsz+mT05NqQ5rCq50A4gG8YGpMe7kBWANOb6SgSnRaaqaIfBiRknF6VU
MNnFMPTMFdfiNdX3s7KAse+IyZObNY81KmgYrwM8avbX6IdPgJafcMsaQsqrNSdxlzJSf8KZGpQT
cV2uT6EOHdK82dQ4vgj+LVEaObFYOHFb1fuNCO8dHT2zwIQb2m4+99TrP/8ja0/hY9SNztr4RoGg
UGZVnpm4/Fr6u4LekfRoNYq35/jugsHHm6wc2DF2jAKrGGdpq+h+bJdJdopMSDGB34udNvlqPGn1
WkFf/KjSp1Jl+Dwgy9po3kSDgkEZN/KtkNQOR5Q6QiP0g54AuvqaUoqpmLJqlFR/yiymWnLkiYWm
tRlj7af+yD0ZdyQwA7pC3U2+RNTD30OvN4hcdPsHPGWjejr3ag8lKZPFoTgVSP6g+gRB508Ed/kh
yVBw/53PhM7R+UnV4PtZengQYxRzx8jpAjEBTCM8mP2Xm1VCVKSUCEORYbKwtOebuDPV6p/junnG
3PJNIKDNNJxGfaylzGa1jTi3KRmVRIw9CXSyP1FxryhZ0/4TxGM/lVo5KQQGqD5jLMoXXOvIbFCq
oXip0a2jBg89bzrVcJX+IfhLdM2EQKpjQFW2AhEWfkJHv1cYn6n0X7dFYrU28SH+2nLKAYcf6UJ6
qPOy+x4HXgugI0Yj3cx2yCQZLcWItfsSTqrFvijRVN5Ap0IetdMbN3aW6OB4QkkbCQSZLaJ16KBs
E5s0yoagd3Snc+ofaBW5/znsgVNq0ymhwq+BvBA6UaYjI3x4BZpUQhAG6iuEv0VwxgirgVkHY5QW
dm3eHMZcdntduRX5BQQIMCOZubS9mLdEFxCSM/EtpDZHizf/QOqS4lFJEQSjKTQ+DMMoOHtS9l+h
MczaiCcXVnefc354s3qA1zBrThzUgIWrDI6zv10heNYXRHZ9w95n6Ay9A1g2rpGd+D6j65gqCYLd
9U/G+R4PamgulSnHxvfednhqKWg8rioMyEW2BcHr1668fGJyfRb2ahRz+V65stiEmd/S/nvQX5ZB
34fF+G9q0zKwzqOtzv3rI8CoJ45zutjSPZn3bXUWEIVwFaqVHfkbXBeZGxIqO3s5h3BF55UzkW1x
QeRqVPnL3k52xk6VHNomETyPeC6VXdxOMLnKilwTKvV8G/63PkMQHWv81l5Uj+hSN1ldMBHHoQwn
7JajhOFF3IAKaHWeN5D2lkNcvcUGPc4eLJXqN9zqljo7KovMxmJztrGPZxvpH5SZ0BFPo6lAMMZM
GL9ajCNyATanbyDNXvZjBsu5hQd2Rv0dELBhkA0c2Bz5GbK2KxYHhi0OkqQHa46BOZHjNldY47OY
vB6QWQpEBlwshCvwxbnJi6l1cYHhSGuPuKGirCdz3eRCxKekzhQwqTArRtIxEwY+hPxuP7qnSu3t
3CKm5g6wLOup4IruC9uvXHA/cr/kKkfWCceNvco4StPKr+PJzADuRwCrWTSCzIJnHUcYytB6JdE7
7nRKDPZvc39ZzHtx49xZ563dQJlioPhK9KTNORP24glFqcuyjZG4dSoVSOgBkT1BSJd0cHU3sog6
/mhM0cC8WLYQi0w2dzzA2T0Mx2UDG9WXl1ZGviIp6kXRe1VmQu86cKHLcKRCDH3G2lt/jR1dCK6V
4uEZwlOMPRVN3f0IjCX9vG1kkJzM8GC4EXPEF6armoqha5BCBt4/qpx0oHXLMxhOlSlp5FWCwezc
7CM6x59j4Cd62M8miWogfCr1qh12cfxG8UMnS4VYNrfTgwr9aTngSBjTaCO/35XXeTusg8NXPCnh
DTg1mSBeQ2mUlXygAk+f7TklHmBp+MW7Cp2Zu5cGUGJ6JYezhWB94F+5QSiKcTW+2zf2zjYlkGOy
BNT4H+EG3ORG8Szaln/Xmt0GP740DTlYy1lgJvJ4RxxvX7O2OLj5KksTET3iRwug+3pBohzRWWs2
Cqz0qVwBAUoAH2MiNXvKcbuJRMlT8b+WMJJxjBvNXVCd/ecpSzBWkUBrQICiAOYQ+2B5WHmK7gZw
SPnLNCmbhZ8Q/mqQM864zPiBLuG9kmlLOD9YrJmLFmQ8d6NMgToqn5VSW6p+8KABnWeFnY0fbCje
SF7OZein4DbHtwlAPNVJDSpRtkp9AuCttL9wdVMkU1AqePnm1/5mILcT1NVNWTDbleZ9CxCHUlp4
avQhGwhvku5v3frG3jtjXnmErVSCQqOqJ8NqtiTd/f5eAv0V2v0s0m0C/MaQUQluGxfTIOeBJhbl
EONaeGfOvQ89TbCaoYMScnqFZevgxPqBYLjzPR+Uf0BjRiF93UWAuTSqv5TPT+bIP+rBi0LSrx7A
PrBGFIkn3xaaFnB0gqf4DgmUACZ/zt4Ssa5OIVAwkbH8X2/BjiBPc64wsPnEoMto/b6HF2PEc2hR
RfafHuhM7QySkTKZ1dtmxdu0uV8o/ZjyIrapzJualBDdn2tZscodLr8LRKkW142GIu1mR/qB+OIU
j7sTQHbYd6VkNPkmUV8CqECE3aqDNMI+bGoTYGGiSCg0ZMCznMuF1lsDMM96K5uAb6PciIcGGG1d
GcVRgiGqP5c2X77Rk+h0nrQxao0tsxdwu4X9LyGRATJk+7i4sOgI48xPyfPtxv1gfArbz/rrDGnR
gHE0g6+zeLBQF+HsABes9FqSiQ54VH0mnsOvQwhLgmm51+9DWAFFy5bp6VRTHEiGeq6f9SYsqXRy
dT7DNcvaZ3DSSVR+IdOCs3OsZRHLb9IjGNXOWkTN0IoxcnyQXAPMBWxP2R4lC0Gr+KKl19z38D/e
2ELcFINWKCpt1NRXQThf7MJ1P+5gowEvkClBfKNcGrZxKxIG+fJ/+lEB7+sONwlcffYqLNIRCVSJ
R+VpdvjfnG/r53dx7Yz0QR8t+HntZ3ScIYfD9l2q7e4kNzadXynBVTF+7pSJWYz3JdEMYiOxDaPL
pRBoIII5PliKHPPoEGxRf5/lXOtXZeFMWessXNHkvqCJD4kiKtPk2rZSJmhZeibt+rloCsXFlwyx
sBh6TR3VbrGobvCGN8Yb8wXRUd04loZYWfmgB2Vew1itGgV9wQJfmmracgz808EvpElU6cXh5CPn
iN46Ig4DW3tkq/T1M++Uy0p5sKwQMPunfPGSURnJj8tJupoutjMeWTYgLIGzMXblBWk7LVKmYW37
YGAoVEYLT7mpxLgenuLTZ8MNwmlT0xriOl4kpvy5py97cNxXzrHtGbSp/Eql7rFxR2T3iPe+pED6
UJvJTa0kJBlCVOk7NWSLX5w8pqak8jiJ+2grbCw0JAn64CB9yqEp41CX/q56VMcHU/NUoZFdGu/M
iBPkJL0/QawyUXvnvSNyR3ErN9KymBNPF6Ig9y987EOljubdLk64lb/2GHqW8ZtA/XRYuC8s0VAk
hsgXAHVPaD1NG9CBxhFkXpFWmsLJiGA7Rf2jsIcZMvayZKGgR2Cujiz2jJ6HIGZqzCeizGNKesIM
B4bHzdZb0eeJQk6xPTWlmZ4TcZ+ZpUHgxrnRQ+4eTFwJUyfTIggjAm2R3qtM5d1sl0AVBn7oNWKM
yc5ju7Ea2UqxSodX0UU3ENLJUz8HQ+o6RpMp0fNP5EDXzBJOJfty1Qi840mV9+WosLbpiFhhiAnN
Ez4bC2nTeqdiWSZy+jRxOmXHJyf/hv3R5KcSGut41TBThImTeq/iiOHUdlfTKCbylel+/cAbUtoz
we05JOSGVcSQOGe/8NO9mhMbXu/AYVOMw9AH0amawnkwfOu2DB63K6SHdvkwwnr1IjL0VsGmoSpD
TrS1UPolidMrdCMhYzGht4uA1eTunxojDUojGSupYIfhWEYwhLpndOb09gzKGnDRkDzB1rFGENA7
OeU33UGvCq2MCzKg2Q8tMx49Ty478tnqX0dKvguDmOhb8BPQ80l9K3guIkFiAje65Tc6CDASHNSO
yo9oZYvjCUNW336X2MyIytM+oMKMsrTk2pVbwlfXxj+Ux5AoaGqt1NOxSjlSGKyD4oQYFrb0JeKj
XfsS51CrQ39ktb0M9preGfK0lqs2oTHiAPJTxvIt9dYwhKLWu//TIRXt+lb87qjzYb3b0JKEoXQ/
U9WDiWLIjpXDbb4g0V3dMcnxRNCPUhVwPMFfr2bdFmBb7OIF1bDbKF9ybzVGUQme0t9wSTpHpWVN
F94DMiJrxAdoINze6CAgnfSszTV+4dSMsPT1Z4GQG1JuWw0Au97nF/Ryx411yjqWNEo/C0UN30J5
mepkAuiMNAk3sNfX3X4fkHG7O7U19VCcnJegtngcR4SIaAnht3RdCtKgyh6xZ++HH7b3w2mHTr7w
DV2KqMLfOq2Axgr/Su1toHvrkVoojojutxO34ZV65wSyDTMDMZqEe6jqQrRgFNSlioAwO1MiCXcC
WXULThPxF+d90zsHwX2sAXe4PQ31O05STz5DiVyGZBvVJ7QDaBWBy7+lSWFUGXp7gPTS24FfvpmE
ACkrZycJtD6+DerCqobEaIhep4FehEdOMryrjmEtV7fBUjPZozBrg/5K8WYGgCrbiHrRK3I3bJSV
DRIhHtBlyg/nSNPSbZKElnM0XKsQuAfqU+5JF7A6sJGalU0WrqBIYarTBnOnoZbkEQ6e0M4A+EvZ
S5Hxs8GEMM9oDIgwsAJ/uFDOYmLx47V91N3ER1gdJGp3f1wDIzC9l31HcJzrp0MuZs4RJ7m45RjP
GIYAs4+lcn0WTXCd0iIO+5rafM2OWq+TSP4rLphiJa/73edN8ffEjdapCdRXFgKfA0LLkYAiIhX0
6ET+gwJvRezf8d2C2mSbdjpzs/BGzEYgF4BioKTYms/yEbiLIR9kkYtXY0mEgzmEfWoxdbgmSCt+
qJbI0j8l+9Jx+kyv7NvjAxJvb6YzL04QdiYqsbLHPM1vb4Ck3Skc2bxVUCOAq2Fp4MiXGlWL81sQ
/92hk6vW+cpunajdb+URnkDaUr0gqxLKLwBKGghhM10sFes3aN2aYci4k2qDduKty4ta45ZVtzoA
2m7Q7RFjhwYi8f2RmwKVg1Y93UwQKLWmfNUIcOPxziP9lFMKyUCxBsIVRb99YlRII54yvrxLwgnA
2fH2wJRVTh2Ep0mx3L+TLMs8/wO/BRqa/m6frmjCOsP/HKLHXa9zW48k8I/zRF2Mbv0qgf3WkP/O
bDU3tCedIU5yuxWeHj3dUM34xoluY2xi8tYu18vbTIkJ8/uXoJcJ3dDu0O8eMMxL8D94x7IIkP9l
GzRo5quk67MhND11ZqQiMBqaia7zdyQhPNVXqacFFQhX2/iQchWrMVM+4pY98r87XUjbCrUFTPMT
ZV/eQ+PZcw8V0ie5SsIjEzBYB+JmiuFBFr7u2WGFf11ZEtv04xZJP+G7s+11WHngK3u6CO0ZuP+6
Lz9B5oNQCNxf0ZvDFxJdCDW7XTpSwNJmAWW+Vk+fRwIZCSt4M/OtcGT0pF8EXUuemSwEZfsC4FKx
q8FWUUq6+s1t3pgm7WHHFHognRIUBGrc4cHBdiTrxE880TjKb0CA4KUmUHsCqOcq15ni1Ct0knUc
Qnjuyk3MQmnsY+F4LjNoGAC9/j5k2BBJT0mHGEF97HIbxQIm2pyFQfz7aaDtufGYqKKux04Aw4Tz
naO1Jh390oJa5HBcG33/rD5mklkA5w0EmMEzwNteAp0qWaWXDXloyDHxex6Kyt7rOq3IT2KGtXUv
HIYgbfMfxmk6C+wOMJJgnzOPvSSxIkBLlI3twj5zjNEKZbPX1HOsfGtpzsdKOpS/tdKN9sYNvvaz
X7YKvoVuAkvElys26PB7PlhHgqeu9Hl8QuYIgBcCSlu/EpalMEsFmnumkuqN/+W46PwX6vNnbEDF
SXf3Hr8NgihtkiD9yeE8G7H/zRk1wkLfsxOze3HkgrwL7Z36y1yOuzf/opMge+xvkenK6YmGSgNQ
ReywXyIIh3Aw/nR5g61DrFcOzXyScr7wy1ohD6g7Sq5rnlS+G/Go2aTOobieShmcwECaqHvVItEH
a3TUq00FN+OUX++E0ORCNl1wtgag6Y7WbtxEhY6lsjK53j25FTINF2CR9ep9rpqBPyFqF2wtlyGq
/oQq161vLWe//a8hCR/8Zc3KjB0XycxS9b6y1bvIwkgIiiY7GFAUbnMPWo8yTz1pR99wHdPPdIJa
xRnzvwEVwMyW/TefngowbvHMFHivM0OuCw9N8kW4/7ZdLsISI8bnsQ2fGM6fjh5URUAZKdN6AUDS
lUGr+tIMZ6YY0Xs17ce3T3mnLlpb6dDjtu5rcDsxfqr4ciK8vlpuj9KCBTtJYSaHRe6oTV0j/w9V
xeZlSQNbhRqLgo+SGmxg8pPelb1MQXWyKM6BGJioY5rwVLlrBI1TL2sTLl4MOlJu4xt0bzF1hBJ/
9GuSdj2nLsUfWEMJLHII5QjhYAuNyx6z4WPZz6fFo6bzosVMOSDUqQfbj/5qi0nSPNpBRxxc67bL
/tMu5F1ObJ8zCZKLWAC2IvYe8Zzg28LmkMT3LKRpmSQ9MRwosntSEaRotikZ+ccm7LOebOcFoVHM
oOC0aSp8m4WiOHu9yggB846v8qdCzPtJaJJ4w0njY5ugmWg3I0JrPc4JhLk2N0/WMstPiejTqRkA
KQJ2xrUJb0Pgj71OsiT5lIbOC41Ez/cca9CHCO0y2dHlArN1NYZwsJ4ApzjQ5RFZfmQoeSs7bR0z
+pb5HT3mtVJyk2JOUPSFg7jTnmcBNIN8ADI+JJhiApVE19tCXKVSD7PLagQFBpdWhT3xyBpf3ZEo
LYCntsQvHSA3DxUf2JPHJOr+7cJcqjKep85ouuypsf1qmVUrezAy+pi/DyQUuq1YiaOitOoY41cH
o5sht1ezdMJULcwwx6r4qQi/y1H45MQsUaG68DZu0nYki8aZHzASAoIHqNoPhtqXAHQZ0/+kLNUN
kDg0AcH/Vu/4Cdurj3pPB5X4wG0wfunkUQdvNQpj4820XEL3OUHZQfXtxl8iUmegb0W33DH+GquU
n0X3tjQZG81t3puOV7CAS6uXJ480DEmCqKN+SblossXumcQH1WPnVW6YjycP1JTPFTNtaWRAU2ha
pExqsfQeyN77xtrisxoYX4n2Bgkzciw2MPrAasW4wjKqYQWnAU0VLw0X3Cd9w1hU5E7HetXsY+P1
1zHgzyGQn6cMb5klkb7R8Q3wwIyEkBnENeDF0Erx8KzhTynvCRMtgl0e7SCo5Rck33hTap4mL7hp
1WAZzgRwkkXzibn9AZBpqMyJKgBhWhR3J9lQKkuOYVQDplySi/COLHfctdj4xlwP5YhvicAgLpHh
aSXgqxLqCCXbAKVtPxjkpEw980+7RRjlAWJIvA83czi1WARQsvmKKMe4HrjFyoRCK3jfEcsAMzHO
jzh9QjnWEJkRvOBsBkJMrXe9R+d4PwSuDwj/G+6Md/22p0ztQjAORoNa6qgobMcDw3puIOmAXZlT
GGSNjAlM0JiCXx7xw0ZjZPtTLJ2FKBRDKaADx0lCoD+emaeg5Qik3q7of/6Kw1yxAZAJXc29hwAW
2OIzpw7XrqNXdrFe+mXvsPiUYWK/GFrKfgUPYACDZa2k1w9unSrSZrI9kJ1cTCS+hgSzHhz8yq1I
0qq0jzLBXpCSfmJMrIpZ7zdR4uddj6LeioLaFOMs4MxEWkXJP0UJq5awkUU8GwmRjxopulvY6HU7
sYXmXHHIktwK2gGvKTqQ/djreJMV/isVBA0yHzk70r0EZkZpj+pBKCM038OMVD1JvFoEl8A5QiP7
hzR+XDZ5pdIUmuVPgKrtb6DFTWYHiMIbzVaLFlC66tvjSCEl3XORjRsyTtYldMXqx+nePCiCwDl6
e1EQVH+skIAjBLv4x+KxuhF/xRwz1PDD+Pjmv/y8cYG7iCfzDoGLvK7EWqDiwMz/lDsig8o+dSCy
NGpb4VMh/rrzxsjuDsf9VaZxGDXWOZVvektJIwqndFL/GX25mPvCOors7RwH7ZqaT4YReoPbMWNu
jRuDMIt+MIKk4CBSYl58o756p9Vc2nWy8HiOQLvnu9HykB7nh9AMo57g9JGP/JrroY86Bo6yURQI
2+o+xkBUGhvfJEXQ3yWYYeflxbQDry2YmSPbXa6u0f2H5E4d/0yd4qaQsRKPCqRv+bakbV/IgcFZ
RnNHdttbBhlLjFEDXuHQu1WVz22C3TN8hxaKo/2U4NJ9WelkNaQQFvHIofVE7Z0/7lxwGooLO8Ny
dQdgJUe8pFe8WM3gKo5lzeakESa0s+5dt6n2ixgRqdkuOzldNpUJ4gCKFgmrhymD9AMELY5R+YSL
3Kgy5BwzaLBe+W1jY3CRy1fgVwKEXeBPntKuMGPOHNOzOb+JrAgZ3KuG2OFk1H0k3swNrY7JWDXp
z8tspu19s+yh8BFqyrVAQE4gzfWVZqmvizrT136vRYaNYNKYFwpLbvYD3Ny48/hEEOPUumKoB6nD
vUZcncRHS2XxcWeh+iuv0N8XaZuHIpaxkWvV94XNJ0kFvJQTJ7tHkYeEaHWsft8g7x0gFw9rrPkC
FLvBahFxND1cRcciQhRX3yyizKIuT+UaLWVqy7SjMZn3/ZG03LU3DM6PBdy2Fa+KgQKQRuP5LSL8
DAewmO5R1XzU1VpiubF+ceEA2e9iw5DoGLt+/f58wJaLGFqtl1El7XHSHzr50irbxRqO0uj5D4vZ
EEAaTTg9mTzoMebad19K+jtKG6ECZNUdbj+N9Z9Et++zQo90RWz9KztlurrTSBuDh9st0wMb7X7v
aRPAMC3MHJUdXPRgPJb9zGzkzMgOgHe/GaxyyxPOXfzJgHlpDtbV8rFcEX9ccX6i3eoDJwRkGx2l
7Zc4N+4B3bi8QONZeKf919XK2HuLYLywZFwm8cemxRJNZotdefOH3h6fc49DxwpW7BR5fb01CPTj
yVnXcZfnqdRGN4MZuKeCYKaD3Bm5N7tHnJYU78UFhSNzUNcsVQ+QhHV1qjsGPVjnnS1V3GWpnJYY
iu44K7kmcvtQdP1k/T5nK9zt1BTU8XlRXfjeVoAhr7PhG+6tw+zHePMlXxL/8mj7syYazBQW5mxz
842SRa1ahkitVMr0X7iWeVQnwHkTHuYBnEybm20uMC3ll3JxC1zGjpvi67wBWzX25chRRzTH4P3h
h2rEOsePEShFpvu25DStJMbxKuaTLyCuXXKCoKu179XuhlaK+dh3KCVk4tTcYzySJ0i9OgLpUSBP
O4zVt5w9y9lir/x3FLAWmMLcgDjXILPMLK1mKoCGu7ZdXcIQ6++qCzt4hPXNBDrBlDQs0Z/uEtv+
2r6tEf4i5ju7e9X4JaDuhLtP8ZSk21WZZauskbZLi3ysjJOKQligCFN6QVY/sBSfxv07mo7L8FtK
5M22s5wQtYZFdbdJQqXeOCTTT8rUhBt6aQ4NhHYX422cJ9P9jl1e//TxPuEieBwlA6USqizuB8zs
EbcARnwA/yrOmSK9R6nIMU1z6Hgff6F0ixI7EbBw85+wk0Yz8cLsvMBy0PkT+Ocm6F5iQk0QesBy
855q4ciD1xVig8KEJ9wfVYBW2Lcrj01V5aWBBZ2kkXLkNdbGKDapBEV8puBaIFfKl/pkSki6Fj3o
tqmIvCwSW23WPl0iRJ+YgddUA2KjYr3E6wwV2UrqAKIkkffRuGDuwYB/6lUlGr0YTCRML57MzJxo
Z2QVhm9SSOBndcvtspuyhj7TI2/aVXK2qk3BH7wuJag94Xz/5ekpD7fZuoCHigeadvBeQVJPa0N6
o13f/H3zNfzW5WkPli+H8Xu4ER5uEK3ed66epzughn/W87cP0G2640MwntNTFUiphEk9mGxO6h1U
+4a/nyufS5drG6cZkoHCJqJTfXO3wc2v/uDOHiRxk7UnQXTv4rjcY2MHFv//FYQRqlP5fsBFJgeR
NzEhhI55yqQUlTTb5WJSOpL0dL4PgCIhCUgz2dlj3GcIL6YEJFnTeCyLgloQbWNH6Y6vUUjUXqDQ
5RIJOxIxIyUtshtRObXYGtgZzebXD3NI6yw7qxs6/Yvqo5NL8cy7Xud57V713LA7iX6OAyrGdKcu
TIh/0ZrxrnoFg2hbPGkEy4bK3sefsWLj9qmW6E50T4+fvFYSs44tsEoCK4qDYnY9emZiHYQOfJSW
clICXYVEC/ShOVp3u1jpLgv3oTljTotzqAf7GyvWiex2U2oIbZql/HpqPpZJs1TQuMSeWlFdPV+9
0GRN1t7bVx/ody7548+uP9VvOaTdU62EtM4Svmc2/4N+RNC176bt3ZyiTRsq8t33fErvZukRpkMi
V2cTY8TcXMFHVti1LdOcFnTtzLwTO+VwVaRnm2s/pfCYO77BW9GPubdwndZZi2Z2ezz+oWtWu+eJ
mMfpUbHsyiN+19dR1ec/+n1ytIQfj3Z6fF06IUYBzKKkDgNvkUXfNGHzg3Nu0vLo4da4OpIVGolM
jwvjv2IDB2jHLXLPxfv1Ce6bnC9nPJS+mo/Cm7BnrzZRNPdRTp1WjJvImzcpjluBWwsQdfnFYVqC
udI5T/CGPSQg8f7U79RClgsWdtdsr/dTYMjTcCMY4aS4EJU4sOGLKNoN9rivq4QRqCxGhTS1Vnrw
fezrgRm1MQaVP9yNwdDh3XUGSsf2YIdiPqmY3y1cX5DXbsQ++yoOJqL0ZBQ8VAZ7ChtJxjLMbNHY
qJUCdc4F3ARbjktC83ddyeLbxty2X6xOwSq09FYvtN8Ye7Rl3Ez5NzA9NszWEvIRJ53reHBfMGIL
FWRvQdje1th5GyXT64y5jvpORti3J1+nR1fSwzrWi1jPKlukU3LGS2tc7wK5Mn65U7LNuPo2/3h/
By5E9HRibXqCA1RpJUXyTGNoIA38kM+OkdqdA/UrN2GVmYp3FZtxFHsAXYiaFTatiKlXiwoklZQu
Qrtsuz+z0aNCI0CqheYimj6CvQMZMFBvbnxpfWFYR9RPnkM0dzOs5hyDUEih19jA2mmNt0EOdhnb
/bsEZWkOGZT4hAfsSrS733kLfgunWNYIPZ/7Z+f4kVCpEpqZMl9WAI6AUwfTy72EfWNhvAy7VtwN
8QWX+oPHNbNcNk8z/pOrzDYRt7b7UM3nGY/3U7PY7SlB9WMoc3G7BknLAuo947RX3L8kAa4yla6Q
8tXGKne//V1w39Ke9z8Bog9meTfCxlmJYXOR4CGiaEwNH8W7EZQnReha/+UdGR5mFpOIGnbI56xY
ammBzEbDajcpDzZiNRq7djWccZyj7KvUh5hKHPrc42y0zpaWj2B3kLETONs6ks3QPHB6qkMFk/du
vyMkFguPbIB+AYAvltqghcWrLzPMxSs8Q1EYyxbCbYF3i0SrI7D2laV7l+GK2Ox9ZDstAWASt1Ej
s30MmIwA491R88q5YXQK++sMUYOC4MzuEgoN+dNZgW7J8Ma/2N/MeGWzTOpGN/pIU6L3ZgMx0lOX
fYbRPVKrdzDpFXOOpUlrk3MUbZVNb2G6Mo6gp3V8h0Fb9gQpDteODfA34XRFjAPB9JAYvCi+N1ap
5bm4BxAAAYHNNN167GiAvmwa5zfWuJSIZ8oH158SYrKdMKIgb3+vdduJlr1uHo85SxGTNmXyBcbM
hFhzZ0pKQWJve4tTptIoCnvrTzSpnYPhS3Zqb1eSZYDS7vIOa3FshWJbSg8sxZ3+g57qzuBGArfx
V4Xj/RtnSOlnsrHmLNhPuHdXBnB8b2hFTzAPtaxEQCUhR8Gh+k0JsmRuBuYTd99D0BV1hF4T2MfQ
+2l/JM/0ejKRPnwSDpWeMeJHmuTOxTfHweZuqo3Xo3bBxMvUTffdMASKBPCBxQcpR4yUktmGtphR
e0z04rMsaVPW1d1yzH0x84XjqDFLpp/Ne2i/ZXDVAX0T3xoCk7twBmZ8Te4RPrsmjX6zW1yeC9hH
XZAcq9k4z/MWYXv2+XJohcgy9Ybf/oSkH9SqYvlS/OH+lLc71EuT24rBDhUg/z6Q1Uu3WlbKgn+Y
d8NAD3e8kPFqTvMSt5Y64cOG9CLB17pBsVzeHdsKb9SPa/3O72gP0rea533RXIBmBvA2mPBYG1Nq
5bsyFkkzIuf2AI4fZfB4OkU3ng5lfAbZsOcVR5K16/lJvyosYI/1Y82/33XvMafuTcypmQkE4Qjn
vfINxAxBg9WxSPdkH4dpES0dDplhYNDV8zyRmDsAknvg3FP48uQI4kulJ00uoFUYk53JZIacDEHP
YnD/z26gDOe1WSke+/qE9i1B6tgt7oc2ERGIo863Klf04dNwxwvwLbFVrw0mjFOWwkHpxZ/X9OS4
j7+V48qkP2S5Qbf//MYnaRBi2xvLtQNl/s2mNjiDSBI2iREKMxRuOu4hyue6NOjKGeI0Kh0dR9/K
FvVgwHh6hhvVxqONVfMc3SJ55BoXOLUlQaxRw4gEGI7NZJo6jO79BAI44F/UtCyorREpT74ixVOI
bCC6XGOjtGczL2/FXp+2naD6VqIBYdc5OJ7r6Voz4NK1nI5bTIEZT8BMp8qDq6jf+aKYZ5qhE7MH
QxzQbOYN07hEXSR0ypHAnlh3LqY7RY7/NfuPjBVoRQ61d8aQT2g8BqThuruLPID2ptN1BxiXA2DP
MWfLCKo0YnsQlXgc6wdETmOXe+q1tjfkaKBl63BP82YrcNw2hEMwJehdQ7CwZFRBMVQhi6UQ+rhn
HFUwAgKV6C2CGf/+GDUmb6qV7TpZFR/HVH59yhbPrFAWX3xI8/sMRvmggnnVcJp2U3t6059lGuqt
luag5jT7ggT6SSRRSQvjOELTFgLSdhZr2zvoVnyz7TBFPAqqCIegrtsrPEsLrD4AJ/WeatiwpVxu
unML7QBcHTvNyLhkZOpEN5V0c4A832YBjx141VAbGuDSB0AKawhkgZswxpwVaeYsieVltlAKYTRf
/IsULSJizhj5ZVAZMnddx9unYb8iZQARgav9ey2vwLgUm1MrRnagFD/zy9b91WQMaLpn6Tw+wMyR
W6yM9vykfgBk1OW3+nCnxrP+9+NxfoW5FFdN642kWdtsH+uCxH9DD5uiFORYxzRzaHK6eSQibuRj
FakqW5JEjbMhdO8zVLq8+Gw1u7XWdQjBIdyfVmP8ko/NQB7/abOgvlvOdJvk8eL1aEc8AyoTKPZ2
/jCjwvaJYmGv7ujPZv14iPiC/zaegyBQhD6sf4waz0/49RmWT2Oqn01vBRkfqA6kXQWJDXryH4IA
9NlUdyItn1vlyRZEJtFJC4ZtQKaDsgJtzqQxfwQCJBZUsdCPumaX6AclY9b/STzQk3aBie/uyvwt
o/tLfZDHmJhp186w4BZxiqrBABfdIk4P993fdjKxIP2QAcSJqLSA79yZaYUDFpj0D0G3eXhWkMe3
rCGQehGtcZoNey/hUneNAt+N9SyeR7LyFgLxTaqGaqSQW0QkZkqAwT2lEvPk2XuGQmars12fWu3Q
+18VaQl3r6I7lJWXcCwDryl8Lo+8H35kD6VESrWduVaiDVsjSwYENSXO2GbL37a54QGenZJICkHU
LgkNJmRF9ciQH53155JzfT+uIPVirSNtIEL6GChQcc1DivVtVfoxqjKTx1lN0lZnIPGNSFFh5mqD
eSJVl+3G80aavsdjJoKJwtG2YV2BmXEaM3DYWEdpGaqbwPt/b/1YKZo/z/nkcbItj0ZK8Ee/Rd2o
hYoRTE7mYZlGqwQEIE4QmG1bXF60ahLGpsf9sIiXFxz05i5lAcCX0lUlXcRE5hBehgyXav8W9POg
XXwm7cLHEG/xQFsK8KOU4SK9LVqCtKAn998q1bEMaLoA90gRpz9BnaOqaAfAPaCY37jcrE8PARja
as7BJDNflI+SDTZdyH4fKPLgihddiuQ7z527j2KuAj9ozsVsxvGMTjWAptF32hXNjJ1FF9VW2WnC
F0d+WZu7yFaoowGw6G7W2EmsmR1fRkbs/vN/cFQG7ZX885ofTNflqtMudo1GGgIGO+D3eOSUe1CA
vaJ9JM5xKztQ9QD2de3BIsJJZl89QvrRnR4NDbJdh/i/HyYUpMXDH9+REKDqNgqfhs8bHvxyKelu
hJjmFmP+w2AzNDP86bJz1d2SrJscGfJN5Ws7FyZwUAp+V5NcDGHZcgG1yN5q692T5qFjhyqoIjuf
oTX3GefqGhvKROoaQSegIPE+CHLYm6LvQmwuieSo9Fe5vOglzG/jq41+k2rTh9R4wOw4Rle1rdOE
UORhdxhM+KYBOE7jYFG6ydqJPWy3K99dd+lUJI8GM2lZ8R9WDK1oMR6bd+du3++Wrup3YSutvPqw
3FShQH/qeLOkUTGB4dQUjaf07AWyAQF4OVZXxZTSaWfCAiMFCx+7s+8TIjlgJJ9v0CWuuNrb1qmz
L1NIQc/lmDFIix3C2iN0zGQlRxQKYfUBcTEJpSqynjkbr82aAQqzIDxDp8H3G7V702Sy7akYHnJx
SuzE5uchBMsNEPiCWRlYXyvbY6Pys6SrAwtIz62f99bmC0chnpAzXRIK1q4OgoKw59OdEXIRIR4P
ueF9UWtNKDUgTYYWDVQY0Bvg4O6AilMx8A7C0M9qcAooeRsBUBRUcYMG8iX4fm5WcDQ+gd4ASE+g
rGBwfgToWg2rnqU0PqAOjEn7ql6XnvZcGN63iFgv8VuUJl/9+m6utGYpRVGIfvlfRTc+hbFJKlxm
VAFqulVzatyYsL+gS4s5JLlc/NV5nqDy0L6T/ADXJN9CG7aZFTPXI6BiJiM9+3MyRCT4z+2vLg7f
5TCYKbx7XI5jD4cmvqGkgn92fvnbqYOslvEIRu9qp5/4FWTAdNixroNWfrJ1LRsA5tMYGVlB9OKh
/c0+7s7dAIZkxdTyZrze7IAnbvbC9mG4YDEnJt8fr2f9MiTWL9EeIy2Z/wqbipqkYZj1XoseIWKG
JCB/ieegoeWSRg+k1WXY+p99dmBJqtsOWzLp9EjCP2R8Bfgho5LRf5hzvdIuiiC8Do8ZLiuVS4EN
k/1FkPA43MPm9WTS82enMD3SOOA3ertxNsTwbU+SHi0TTpa5/SDi7WLJKJVjMMNxuiGH7OwgD6Ih
S4o9uxbnIuDEsx29ZWzE6sPV+zjjRxjHbUGzVYVxMBtFaDve7aiutMju+e3Miab86PNEqlHYGUK5
WOFmRCAeY9QkLUaxPVCEbTB8mpAd/XKjilg6s/gxjh4wFuYNUijNKcBPau1Oxsakymd8/LDVp8Xh
REoctW5JOgpcs4NTX1L0Fl8+xZ6GBmitOSRS7nSHkxrqVSwNced8mtnUSfV8g2/EoDqxDT44JhEv
knhiWHXv3om+DHZTp8NyMkEOJ6vuhSjhquNxHN70NMdTEL4Dvui8R/KikJgH6wfIMdWPq5tIdR5E
I5tApaD1cd1nAs5gOsD8/c7mt/EmgLzWQ7ssfXmfAdOQyD8HOVd6ECCKZVxUwonKnMkB4il08SbB
gT7pahjfSJbqKbEkJ3QBX8F7OJWhxWn9IytJ7WTGm99TaiQsZeU9cn/E9G8ZgIdtgb6JmMSYKamv
/KqsUYNDcNqCw+eNpSgxxhiAeD/rbQbl6dbqey0Gekdr8uJlpmtg404FbC89Snc4gcwvh/QD8Ovc
NAHHPDSpOXIaRRj+8MMSHWHH9SrgaXMme14d2M8N8M8CRJ8QbFQ8h6pN6vSSnrVCkeqX6btAQwyd
CRt78sxSJITOch5M7XbDcVy0DTv8Av7RFgetupwl30TmBVy80pR9LNYsqmAT4E0R7yPRQUXBkSxL
wtRnYEFYj0zEcAtCLNUVQ7U1PcDmZfYgAyKkgYgdaVfKS7LjJ1pBJm7x6a4a/VAT7S+gLpR7FCPz
whLBDxuJOnx8v+blm1FCQLB+ZHQ/sU3y+Ax1nPFXjaHEZRAqeobr7RUW69GTBGBSkHYLUjt6zObd
7445tL3VUhb9kW7Jen+DzpoV7DUYzqc1M/H8421meAv+ZbLMueY2Y9AouuiCfIQRklqpHQ5WF8Bq
EfbtCT1FacLc8BG8OYUV4/xPKB/jVdTVH7Vp4bhg6s/xvizk3L7G1BMVWQhB2nMasSHQRPuNwEbO
x+0u8LnV4ZZbrEuonUFhysRB4VL0NR8zkaqNcdTEIAz7MaXZUjpFmd+UPwsDDllxDB00D/1/104P
fxX82MkRl5FcK0xdnfkMr2xFGUIY+ZvSuXQKNhy4nE7nEkAtjIPf7G3dLzlpOyHWTa1ZMjxr0AsJ
0QSBL47UdZGDvvGh4dDvQMxuyOVSmPDzkZCpLmLtezVGh9LDfOgL4wFzc4M68o9GzC3yORoc0OvG
w9tS99zuiXbKUba1xtUTrG0utF0Xity6xw1RUS45YpDgqYEUrC+wFCfHsVUXsJuNiPBM+B1pL0qS
A4QgWdMuB9rwkM7VX564jK4hX5MEMYa69ovgGopglt+NbGYWo4EtcCGD0eN2WcUVua5FOCIqof73
fCV/u4RCc2IdFl28Vd+CtzSZbMWqpkfAmAnJEZIvMzBDbJCSXyCBdtNUXOZ9o1vvhjpnLAYDtqsT
RPyPcIlFigQSXpuxL0IQ/A2/Kumh+qZsuOXfjU3+gurP4B/ZJKpYGiXYSxe+m2BvfUZW3IQTEdpk
9bFfjKLpo65wtRC4hOBeb5srcv0GXgrnZSOgqkevzW8d1MYkQwHZB8KL2C3z/yLUEBQwSue5+bps
JTyggzUhnX50PBhy5PR947HVbGOxnquwUdVXbAv5d3NqgRcl0FMemYbMi4DRb7ye5qFxU//jBk+R
oqYG7RQR6qatn+8gh5jJqvW1/9uUoIH6s1GBIlPHuJel5bUy1qG+uwYAukUBJD/26ShqScoInx69
/ymdPHXqAfeXYw0Zz4LcZuCU8dK+qbc0uOiT0Q1LL6GNatu5GXyi6ghkDsihHc72HBYV3sB4Dj5r
vI7v2813/nYdlTktDBws5xoG0nOTs/UNAmuiON2olQYBCw1FHtSWgHoJoiL3CHQMDKOBcLbPuzcE
R+n7tkTfQrYK+b5qUlC4qd9g41E0JsmA+VkND4YWzUuFF47w1Re0UCQd9yaM7qbmQ+SiyDpMWOzc
cYYQFar9DU4C4JEFKntFTFiTIjiLIsGpb5ro3aBuRTAv3zXvGs6KBTV33z8fE2z9u0ZCCC8IyWrG
aOpb/ocqgOA7obDvgG84Bs9bPaAJofAqSHYqr/HEtQV1XtD1pZsgPHj2kHJcEboNGkk/+QIW/5zG
1CUIDhfxB/xUsEcjA9Reu++E+Orq2A/adg485VH0uzoFI3csvBjeCykM/uQBiWeSjq/2wDB3EbZh
Sp++8+NOxhR6tUmnoCBNusUsGomSdR6KeAbCRK8vjZJCeU5ol4bRye+F4ZU142QBpKxJ92bqai+M
kp3pSNIaxyhJaWIuaZzEXGVcHjjAM/bMfBincU4fNE0lpoYc6b6w9rFTuBJdkEWijnTV2Vd0IGaD
nNcv98UTyp0pzsJOu+IgPsdg+Z3jrMJWNw16LZRQ5/dIpGzAy6JkCfWlLaK4v9KA0ZGrin4pZPdY
g8qOJRI/o4PHitArB4OVVtX3FvgJ/xHVICervZJ7v00A8LGd1PoafkTORxRBxXjZp2MUnNkfkrXh
woWfOoyxxJB77fIkELmUPmBGaiqS+JDtuOF8dgPoelPOWwjMWL8vQ1oF/iJ1wxWlFxdMeldUhfND
RtT502buHtZVt6rDZ4hWCYh4GLxKS1RZnlZMTOZcqJpXGE/0yEzc4W1+fHvdLE5PP7k6TqJA2I/M
94JAflh2mQX9cFjkHHie3ef3gT3KXBQft96C8gNxVF0/36ftSRIEl+kZQvaJhk34L/GNsFx/sq1u
bO2xhC+8Px4fKjl4AxYEjB7RT+gWT6QJHgx9U8HwqWW7OyCHjLtlbgD0r3B5++z83erTWdJqfOJf
YHjSfKfGDBB81JeN4iZw6LjLJ1/Tum4v1ayFt943+pols8rwGbHkFr7K+UrqQx9OyULbfthX8o7V
bzBXvKMJHcnnpXIkqLiCXVDLHZUZqYg2ctA8THWGg9gnS2vlEp+3RuKoRsJkWCTCLV5ri8uEniWa
252CHjUvnAcRw4J6YqVu87JMYsEM5CBTdxI+z738HTndXJqx+jYUYieS1kK/M28dTogIKgeGZIqX
ZSCbdZyhCQAr6poxAkAGTXYXzN1fOv8Wzi8GYAUjKptTcR1Gmjdjv5TJgQ6Ytg7XRqHRWC1oBHvy
0NQzbJkwUgm/jD3goNmwR6ATSzLXEubuWWOT8ijMkBF6Du6UGzHqyBT+a278awA8W9SgbAHDvSGi
tTQuC78wRNrnwQxU1WuYjEKrzI16hfwQWrkTQOTWjhnes+X+XJu6xHnmQIG5KeQK4RLLX/TAz9k8
3Vizuo3+cC430Ub4IOYB4Ehmc+mWpgPzk2ALjecMozX3tl7K3QS6w6XBWnH6YIqc9QurCeWM3wtg
Lety9Fbmkn/uT9uW/gaJ+60l6oWVMXpg8PlH+3YMkMK4U56FB7ROF/yJTvLcIRv2eiZe2B9S3Hve
YLzSWh1ev8K1jfyyZQ+TFV4Z8Mx/fgrXCqBrgMcqJFxwkkFKvZtrXzVTceU1qL00lx0Bb2FuTom/
PJdESbsa/DATwPNSIE450l29oSElNKhhrknnVMBVU87p4bmWh+SC6ZlDXBIChhI5fQ2pypr8KKgR
SHzo3K1NByTn9qsB6o1ZtQFsgYnbUx6eNIMrDB9D8DFO1QNzFIodrQhuVJZL9mPcosa9WtQ2AgOn
GgHHx+Y9nqNDBHVGZqKsOef1wDg9/WXhkfm4HA0ZCpE5IotHIQntpH24XUhPWX3XySOswPC7l7fZ
E7pT0vBdtDOIYC2zS2lU2uzVDmx7ow65p/H647LzrNt87nuGSTKkieuRO4IzEBZJaJOFGb245MWh
B6Z7nGPKl6MjAgvPKB0V9PxZ/rBcwYbmVVGtxbT0+NdFQKgjLrKGaIQ+0l9UdK/ZMJu4FJi/RHGM
qHfwE7nv17WZndR8oCsoX2QwnGa85qtJT0cykkMKj4uVjIBoeygtJH54k4h4yp24up0NAs3bgaE7
8fT4qrUE8AsorZ/3M8su+GfJsLGYLTWW2lDbWFI3J65ktFkCld5UZou8wPjd4PK3i6vQaZF4DWv+
HB27PEVPxSDOgiMih8Rd9M+4mt4W8jztoGorkrGwHyLO/Bm6Bu0FI0JW13HbcHbpSuG8VOWnn1y1
5mYVceJ1eFKemhkXjlV390/4QyUEzlm5F1VLIKy9iiTFOjM6dx55cqNqjliv6aidYKLi4aziIKme
m2WSRBBZGkmNMBm4ShPoAHv4BN7zfGKkKBLuLP/1E/d4ctgiN8VjwJiXVbLjfyYhafAKavTZ/Svv
f+U1jmBUpixKTGRA/mYfGvdClFO4dxK4cpt7GqVNKUxbEqbQKMw5rujoBOHz8k83LPaqtFmLBp90
tvYMlJwpw1MFp87MfzyUOOiXKEHlXenvvCG+jlkm8VssbFbPS7AN0vw96aWYwLx54TbH+hEGqlmi
4QnwPsW2QhZMnRvctWppyoyqDdmLWmgZ33JUcfvOF4uoc0fsS2DEQ3IsrZiyZLrpAKnANrHlmw3+
9jURU6O69xEfDTUEfcP0wnU5joi8K+CXn2dzOT1ZFerJpp/1KktKqgRPCz+4B/4savNlNDRDUbsk
NCqnwdeRf7hHcR5yt1IdLbxEVn7UNNAuBa+8ofFQ3/0T89j2BLtN9zVJmh42HuxbTrxm1rZBVAgN
r+yQ/SRp5YOycyYCilQWE2hG2Ex1F8paTr+Gd+6n7y3lGGMT4fTOL1sg5ONcWPjFi+Mt+ZyeYb3t
TadRwD71CwceDAbePqh03MLD25AFL8UhkSiSv4afwubdaw1GKGP0uaFqPkTKyQ38zQZyEGcNOx4I
XcAkV9bBxGsjDJ+yCr8SVjWlOg+84lBLXHv3udZsBvqzefZloPkNEagBUaR/L5dcFM+3M8sgeWw7
VneX0WR3vDzUQx8R9Sy6pUKxw+xGrB0zEymNAbljId90lUYMCfOOoql5VCZuzuswR5VHcCi1YElA
WVAhMbZx+DH52nvljKvjVZZcE8Bkv7Brx6VGVkV8sB8q8zCdlbMW43p58mhRbigMJVfdT6q6YmKi
UBG+Q1bV/toCHKjV7e1kMPqTHfcW4bVh8H0rDCl3BItkmG6t/S3PzUN7IVjVM5EYnHW/ShGMQ4fv
n4ZZ4PTYf7U2YFpVS61kc89TDtyupEf5ehETODpmqz0yYtSLGNLCCNrjzqkPQ3dVezd/xkIW4tXk
FdB3J3UcKYBgBr7jwGv8QHJzT9ExhgxygXtMcOkusDQGnd3TvQqfvOuAeobj936UFd2bb3O2kMvc
R43NoJLRdHNP7EhJF8tzZDm3ckAhQ9DzTp5RWQV803mOpLxgN5ZO2PrrZ0u2mWZbg7RVimKwlZo8
ePsX/UqPONLbG1KoO7Zb/6XDhWDh0xEMO/C+846sXZfswfj1QC2LgQn3rKDgpZg0yus9KDICBv24
Kl5ouu4gMpbJJRFtWvMUo6IYX8kdHn0ImF4pz+z7tj1i7yWa+TrRbDbKXCnVuu+8WcT0KPSf1LZj
/p09JKN5YkTi7d5xzS5GgxI+l5LbUyta/vZq03hQQyWMgYejeew4t33RmxPLUvEMSXIr4BL8wXeT
HfBinhd0ZJdRyKQioja2JDAADwhg6Wi6eOvgOjgu//9IPV3HLQV8t7ebvCuiGJ/kyEFzt1gKBfkc
0uuUARMwO8T14CaWe/GTf7qKZ/pPjN9gPFH6N/mn/nIPYmwLu+3jEFl3z9kTrwI6CdsESjUM5B1T
+ERGtoWWEAz1mCj1ul0WQWcds9DC9L3KFNpRji0Mu/1G/tYgNDdGNnhVG49vXkHk6rv1eWrRWLKx
eqiu3rw4DhTvbvWz7HvJ80QK9AfRr1SAsHFbOFB+jZS7Du8pZ8MMU2NZMk1vNyejT5sTcvYfLIJm
ZB+MT4Kktv5Z5xKlV0xSVpjJv2GMtuPlBRz/67LNVJGQs58BRMKQkd+/vhntQSuDmoxtZInrJgf1
5yBmkRnDb55WkvcnbQv3vvqPuM7kIYdNxRXnB9FFf1mILxMAvXkaY+N9/0hC5adnqjjh7OIuu+B6
12M8GTxlPCTKv4s1+mi9r7W+25mK+X30TeyvFNZhu9IRk7YSetkd4z/UHTShpS4povmhASJ+4J73
CRaEQOPci2qrLxYd6WRTxmf2C20hJs3b/Y/rH8RWLtGoa2xIy1bIrRP0tznNBj1sxzzTH2SM7+of
zHnsSaWK9Pg8LcIRm7R8yerW9QoKHzQTZ0O0hbULhlyAu39JJTwyY0q90rJx8TWrYSliI7ibihpF
BmOeOENVt6/Wlird9i50gg64lyLecXsaqpE+NLUVoBQu4ylEKms//RzUM52JmUTenvS5XKM7T+jT
Z/21Aqe65y2c5uWBB837RKuGuzxfeYZ+agv2/XX56oaZ9DH7YycsJjTxUTmOqjWB3n8w03Y4yGlw
ElC1RWIwKaiXw/a4lgnUgkAvP6eZYzg1o+gEbvbUTxCQ4qKFrkaOBSZOu/Z6AgeQaLiOR+R2rCD7
D7LYVCA+BNECLA8ekMg9vilH5mCB26enXdmEbcsjGFlKEy+dGbB7bVbTbkSn4UzlDmnJCi+4jdf9
MemkrKHQvLtz3m2f2a0PLTTfhSUXt2MJmD9c9o1OIVXFyDsq0bAk2oH2jZ9cpX0RiucPvu66Xhx5
ar5+1eNHGpMwXSKV4G3qx5zHX/QzH2IJFJRDf3d0DhPijiCmVfCDhzgYHhcTjMECFmkGorLISZVg
3cWQ5YPhW6NWEhfTgsngc/gWtTok8auNFzH+7BuRQf8DOoORUZyYRB2+tlLuxfFkJIf5pOuCBXUP
3zGERDaInNspa89ulz2+c2DuZLToHUvMTZo4SxHG/2PXD+cJurzERt5mnvpOJgoolWii6vEK2JB9
ktZPeon5FtXgpCPM2dc/StnVsE69QZQNA4LarjOnXC9SjUNods6TgWERbFJr02RshXxMxeOt5MMA
I/XXnJmpHpgD8qtwR6xtTwD/Jg2FuStEOya/mPrExZEL+j+oAu48NNVLkJPVT3Kqtsl2jWeVzKHE
2PbJ76BpXxVvRKV4g1uyyWlfDt5RW4v6Dur0W0ltPSXIzkIl1Rzy9aNVwAm5fR2wsJgUdicbSb+v
Gxt/DIPksR3fXXNrgK8WSt1L4mkXMGUIGoR06OynF4jv993J2FLrNELaWkshFXuG8eT//ctY616A
j2ObdlxDl3oi/CpPwppJQ42V+ysbdThO+WnRY4WGM5+Nptu262J+6nhE+/u4jHC8yKaw91xjkjCo
4NGFl1xsV4aD1k6BPifzNYTpJPtXWhrVEK68vXfLKakQVS0moSoJR67HIy4pglymt0irOONggzlg
W7uAbhoF2E/8EtGuE07x9q9dewMqESTpCUHxCg5hh7LpC7OEvnHiuqJlm0x+cEyUN7bNqYfesV7z
dk3Tg+uWgzf4MivnVFenMH0A0rBD7iglLMSkr9ZfE6REDsTAoS2eIUzD6TqTLCKoJyVzjg7FZ8RC
1/W6FqhQq2ILDj1Kb7o2riJt99wq+Eow5a8S1v9dpTyLaWneZ8bfsQPaHdvEqTtd9EuyxFBBVHSH
/L8Y5eHPG82ZOLh3Lp3WSZ12mPbfpMuctDJNobFQZc0u5DUPf6THzyLt+QL8nx5MoN7E5mNxbNj2
A4cx0QWjwPW6QaYJ7lcqe8FUrN+ZHzbvmAzqVGSUtJeRLwTbA9SYAK8qitdSRS8PBWAStP+acZOy
bI/Jgn1SMtU0ErqgmZGofom0OfOF7AWa6hFiDgz0PpFczmHlEHUaBV3rgx7iEFqdMteGS3M9Hw66
nv+9DA+nMfBvGVBGA5NU+4k/9jrka0/B/99KrAIGozhIZB/kP/inhiDfTQfZwHAtIw6ACtzEZ5Pv
hDrgpI8krTzZ4pvuyD2LXhVNvCooT2OH6nwWjoV8pw4JfZEwaqiC1lJcrjmeJZ75/h6LZH4cUVdS
XFC5i+iAUUDF8tgpb3quk4Vo8MusnlYYEAvVakpw++gOzs/UkgahJkVXyRsZSGRsKjoI+Ly5jFeK
pYf1EAt0HUulaf7whuda4vmtb9TOHu+/vXCmO/+2O9S7FP5cqF2Hf8xmP7yiZjSL5bsl3UExusUJ
j2lJWaBba0HtBZBQrBRbVE1E6NDgim1YgRybxtgQL7EWIXcJqavqM4XtTJqOt9jj391MKLOFZOcU
JLU7fMt30ixuX6Weoid6aPFdpsBWdV9o4ODKSifJFSPGGW11YrDbCAR+Y6esEG1pHr9r2h/JLhEN
mkAL/3vLVHxvs9prdFi5Z9ILaMn2AOg6yARsBSSrDFbR3rIScFxnwCT4CWMv4suYufYR5WsOdWg7
4UY+U0R+tZH1QShCx0bPTg2CLg9MUZkdDsq7/gTUVBrf3rPM1CNCf5F/DeM8+mKIl+EEr9BfW50o
azQE4TAhYwtsEBn/5Uqb/5NW5mt/4zzQRBhrQS7ZYa7+aM3na5Tzc2GqZF2zhG/L6CExj/wUCHbz
1B69cD6NNvQYEB67NmfGFOZzP2f4hft50UBOWsmK1VH++Tp5MAfwK9SPlKrhJYoMnmSjZhCPHRZn
GdUGAeMT1z8LCPeSxbHc4eai2eoKlkwQQEYCL4n4YSM/JGshN1pZhaSsi2368rgB7ytvA7QYZzcX
ZuyvtgsUDMOje0fAls+7xiY4CX7bz3/hKDqzrp6wv9T3hDLCjr21Y6YwBKaE+wtZVgG8Z6M5VM3e
6TCSQogMzVEl5N+nqJl5hnjI/3W0/kC7374HfSFZncQDd9NoU8N0uyw9e5SqKYhIyVokOJeLiSJM
qeFTNDygeGavmN2lo42egkrRWevg+9Xe1lYKKWOuj6TyUaHK7WRIrLTS1RPbR612i0brK9lvvU6T
y7yWg+84MEtJ2IhiE6I5aAZRvYzRFIF/kinGfPM/fDZVb0QDUw5dIp7Y3RQPv/PUDkX2VodDCmGV
Hf3lsmp0uLozM/jA+OpiUlJa4jMlbLhr0KBpqlF7ZR8wmlbPooDNwLm2XHFwvY9joz9CXmwv9/eH
dcDGpT8f1kmCBY+FUSx8qzf2VlXACoCC2LCBeA9gYTLb5EWChtcYAi2TuKVYHPMHUamZBsBXWCU/
1q4yVT2XNGrZp9MMZBpE5RscuK65i9If9ejbgWDt3D82bWMYaO5n07NLfQFQiiMPcEjgQyuttDLG
RWjJLjrFKLpevGSY+TMiP0fva+2aa6c/5E4fYJK2MjaqsphUjVOMj8ivmX2fuEOr3FAhY6vTBsBU
n7tUGesZBdLWJb/vjNad4KM58OyF7Zxrc9DSesAqLxCSqJCj48pyG9TYhL/iEwDfMttJvAM5TxFi
X5YOYyj/Qcsg7+AVl9wuC2hnvCO0gvx/BLtJZK+hFo2h5dHblk1XJ7HztTuGy06lxQ90bVqg0EQ6
GMVjbvqjvFA4doGfJ2JxfA/p6vejev4Uk7fUhqQNG5/5gO//HJilyV95brywIji8pu5DA/pv0WQm
aZ3g89BCsgAI6VK4fqFFiJZPBvDTud2/BnEt5Pd5Bb3uLYIC5CFr4uEsXlpfuZZDArdtHx664In6
skLriALeJ1Ei5TF05iB7jpWE6WwAsjPK20Co7l27kaPEkQSiFPrMvJNrZPLO3/SSA2XtbVbDPPYo
fDc9wugg9qvrHEu2e05D1GnZJnsIVkwJIMEYyS1cUx5O2qHhSQBLnXOOf7RLeshl8xS4nxRiGvVs
zAkmK3CaWsIdyCSxXYlYg7rl5FvyT4Ho62lLWD9FNYKydXBZRBaJRIN8MJ1NLm5wlBsUO7XjNVqP
TEmRER0FfwcIm2md0jENOtZAzpXWZVfvXXnhgUrGM/cVkWLOJyQ6z30enlfjR5X+9MrnDdj8cLtQ
Cydmd9G5lxcSdCUQviX0on5UIzl41WntZe2RNT/0AHW7Frx3RJRloPT4shw/IM2cO4tq+BAW5qty
OatmZUeOyey6tN+5jTJZs1yuN+unPt7XbK7/TAC+dd35dzJo22MMVb+mhTDnFiwGblXlFmAjV3Ma
/43rMjjFJh1gs2n8GgTwECf8n1wBs3VnRHxSGxTXsf6JHAR89rmv1d62NPvi876y8rfrKMqaLZhR
tCgZ7FxMFXBj/a2fu6jjtyEamIlb9kquwyi+Vs2EDPbLDyAPN1uyyaxIJ85RLCIRmr8g8EAGXCSA
mR+kEm0FiZrXmYXOkoYaru0jtlKDucbUWaDvoq3DII4iaKCZ2DGBVtRs9M+befAoQSC14ZfoAyVr
IPnmswZU7Xja12guRGbkQmUEufY5eUKeHNZMRWaIgtkoFeH5yOvnGkpYjKpAOp+rVib/9mqk+Is/
zT+z/AVjrhnx5m8d8PjgKhd1ChvkB6wrQVc7R8ijBId4zyDrm3eB8vZT14Z65kl14EXDcxCH8OkM
gQfFiDy5TfxsxrqotFZ4nHVlTDZOMCVAq+XNQFxT1te8X39BZ0Zk1BfrDwkN6LRR9ojLaAykCbSQ
clv874QgtAaq7qaZ7j3j+H78xjnzHlKbxygzSHj0xiOjNEhwbzZ7Z5C52ITzydq7fQdsa0pePEnf
LRV+xXavoyvSIoGnnD5ucSnz3hEl8w8a+DyJ/QSAts/9FWNFODdYWuUdk2dq7shEPEDd31Sqn4Mn
r7e/WnU9p2ebyI7ZQvHluLrpAaDdGNCNyqvHrIolNkVl20Jx89HMuauZ2YiJAQRJ4MfTP584xhE5
qvpsEt+fPk5juGBvlp5g98anwAF2XLVpkq5e3k6DI/Ozl64VrzmYHtcdzoSYcUmrr2YxfszAXrnP
2RptFSjG2Xo+D4bH2O4J2b5jDwZ+pcnfysnf7yFu2jk+rV16i0fTpwXVNQo0z4ip4WzFN9tIWdTG
wsMuka9ZiBcuXLYxFFnUU0RLmkNz5sRgY94daaCdCV1L4bLL0s9VBOKosFTEQ4gGLTpllH4fH0gE
KGFUYR+clZ6FseYa+zu5rSyc2lqVcO2XGHPLxtrvbV6YdKwO1ePcjpbd4yAvS72Gc2p9pOijv/5h
weuz40ZScmLnJRE0m2krHpwTojfsvj0rL+wSMYYmmf7TsQRVphHQbejXp/0SeaRDKbO1JlBxJmCG
7b7yJtHTDyKHJm7yvgOzzyM2YCt6QqaOHqG0mALmqmBJUkBZvYS9Hgx7Z6Rz7+eaewWWJOC+/s5O
BIxCVICqkILSnKtFwjaw8zY1fdx6v6Xa+pQmxKnpEaLtDhdoJrhXRXyJdxPvQXK7BbHNJ1nnzsIx
VPfOsyBuWnspeu/2FAcJT6HTwMfnT/K7X/ZZmO/xhCPPBFQn88fjYKXO6lfjb/G6pGvR3Xm6oFXx
1pVsDqJuNi2EFZGzKlAAUxcXrqW5xm/E//pYODqXihFsUMxZ7xzXqhA14q38iuv5SJWUCdVoGgxM
IemWCmbpjVFT5EP6ZL+huGzFSCTH4G0mn4l0CxL63EgEE+hIX0ArmM0Mzl7un5uD1LvyUSTJ/PPR
wLmZfbS/pQeqOGFVb4ql1M+UTwtga9x/Jeu5FqhTGdwk/zWKKIQJeZc8iqvkSqOcBwiBuuY4nG9j
1ryRTqBsMpJz55SHbJB6lgBUMdqlWghLzJwpViXv5CoYPM/oM38tvUxkPceFXwVe4M5tGPVO1Q9m
TvoFPG1FZXwy7YrsDsG5ciTGpj2ht445D2fvYMg+eMHPIcwrLfFlQDRdQDRBedQXtjI1phqU68kP
t/firpVNiu9d1kiTRZsX2gnJZGRCjThj4rHzBlCTJM4Kfty2lVfVS/Rb5Cg8KSk+wYci501Dyk2e
vFgOQxFN9BPOqEXAObo/Vtp45jcG5KXg1VZxjUalUJ4cNVk5XmGbSqRvumiOI2oYFuVs064x3i8I
n+FMYMNp2vu5JIcoD5Cvwi8Qzee9s8Sk0CDhux2qrU93XuHK+pwu4Huv0kfim4OQCyBYr86cPExp
4nQieW0ikGvvxon11tkzpSAdZo5/pH3BaVSw+N3pS7HX+Y71UN96A2uLdScITwvZIucoc4stdDpW
KKsw0XPDjbykiyzIm9uCo1SjWBdxgOD7WsoUjxlh/gLoMIODmT9bk9KlVnRG0Va5EVibYR7FeiMd
w0uypwIQUF3AXcf5ae7Bvx4zGEpGqbn3pvnnfK7zBMXYGBkfH8hau5GKyeVca5JnzjvqJ5HKZWdP
BpSQKs35ujSxQfCxvJ2oZmAQXcZnRzz4PIcUT11PmhObxgi9Wm3BdFg28eH3vi82rzzb29iBEb9Z
KR1AqkSgEaF5QRljd32Rqx1EsRgKQWJZUJUiNnvJuyWEIKvDSZhH/lYrMTJT5voI7l4q7q1xXr0H
ggdgzFKEdPSIIffoBLpdtektNlSz0Ecl8Q+9ALepJiPr1FBjX4BliyK83TsL/9Z2uamkryE+lQJC
4xJaQMQEH2A6EacnNUeDW/OPv1DAYV+zj07zNARu20mUZFU9M6yMMptQKHeSmbfZI9AXsuebQB1J
1FzBq9KTApVvJyp9bYOpzb0+frszUVh9b2CfG3D9P7dGnbNddOik81KIIUBTkvGGkx0mfOc4X74d
wvZODReGkcXud2VKoug/lf95JUX72iTUmMPcXOUtCF/KYTci3oqYn1uUPXADyjqLFKN+pwzOHrWk
aQqu4Xwm7p8lEL/cchaHje1KP7qtNWkhiBgsFAlKvsn7mRBKAhQLDsY8iyoIxg5Kr+tQ9VMn+1pJ
3LQCDo79i2+WiO9gpW4pAZw0yVFLjM82iXap0KfjdTYeYLptyCDf1R2aPKAzNG4ra0eS+fwtfiom
Y6jRro7WuwlAwtknAfLUdspyHjZR2btpm/HpFW0ETAtseMOsLIAcfC8RAJIYv2dlXGV83eVSxwcB
vqXYmorO2lzx4ao5Tu7W33OLK3/hSvQT4Ny2iL6d8lHE1D7lq4XF/FtmnrDRs+b5EkjD0d6RM6a/
jSPJhzTRUo1bUXCt04LuLJHeWV5VN6ZQImFqcUeoxdLsk44PX8duvnXiqCO4OUrQcjX3E0zzl6y2
vXNmNRlPsPvg20g8aUjmDvqjhI5bGJtQA1IG8TVr3EJIuSOcE2nba/xwnrI6QjDO0q08vkIdfqY2
xrf3YX5kspZsBtl4rT6RnniKnMKBsTL/9teKD/3PShiUBSx7AePaa13Lowool6ReUyWu4qGimFs4
W0y3Q/bcms8Wdd+NEvmgcPqEoCr7VHxWoTeYUv07eBxUzKaPVRajjuiKI5Pet8W0wewkMk175Qyt
m+mSJxjzOqRMSgGLX7x2RjZXGykYzPrkOgAKZ3daiPWfRLRz9iDcIEKySJfojg8dNlizdCSnCmgN
MkLCLDqoOhvUmCAMCT8SGy3gdNl1afQgDeulqtxjXPrGieSZJVNzFWnMde3ykre24vtxH57y/7Tg
+7q17Oi8XxQiQiuPIUUpPknhYIUYhZvsAH7w4g7ofqAOHWUUEKLPeCs9h2GQrTO+aPbnP/XaL7hl
2dxcx+C0c8tMq3k5l4J0WTvAJVkTquC9dEvloV68ZNaUMzDmmozhab6LVcHJOUTe1rnVSq4LdDeb
PDOKcrhew3U+ZFkKYaCaiOaAi9XBFwuWPH40HtXEtiWqGgoEbJA5F1VNgxBf18l2IEalhMXO68f5
5+FSFZRw/Po2hfdcBgC6qS8W5hh58zo1Jb9HWtY2x5Spri5muUL0P4PMKUhcfpjdQhUN2jJFW8/x
zYrnYi9G4p+iJaXbN8fDNII+gmR20F1jY34qXfEKAzy/U/p7S+OHn9HXT1xeuXxQLVKnQx7wZB7e
0sGt8TS3N21bwnNADafXxaJauh4paT4Vc6rDtuDtPN9YQJJdcSLx4CFn8j0rSFnPbS4hHawBGdzC
ri87qxFEaIaieyZBnn+fV6GJRskw5StGlDOIVZLHMYeQWL9Omm+pQDB7PBxYVPsZYUaKTUHOnQBa
73JEeMmgFg4rqYNNy3LqgmsRJeGoancxQOEYCCpulQXIjcABrdWYTysz7HSkkk36c6iIG803g4+6
YwFaBRBkSy5501SRyjSpz4S8JKe6cX8ZmD1ZYEsE2Sq8e46kmCdkzIa0TA++uzn1Zd3yoEGqZ4d3
yVwzp49EvsenbJGOL/3K8ueKWZ4Wx8XqPpSLyG6bdgvxo8Fwoutt+vBUL0iBCdVrowLOaSYmvdaR
cYUBfjgI+39ex+tutVsLfEq2Oiq7aYS54p9hC0ecJ1aZtaGOABoyoXj1xl7hIBKVqmDF4JTGGvTU
UFAnsBiRj4izNXlr6wgs+Z8m6nJJzDn3jgU/nRbqlOKtOUfA2FcbH9sVT2yXC6lYBm9JYm4vdHXj
FzHJUoo6NWl4XTYNfhbDCbmHq9vJnVZqJy177W1gwU6I7b8U3DwS02hI9lL94r9abvV5M3mRmECa
lyl4NAQ9tb/a7Q3Xxu+bNikCCGhEI22t1DiEoflgzjzf8KdBkJCaxNUN7EmanOsFyaYHl5HJjqp5
cMf7YBOpCetCIkRThmqHyCGYxfpYO3PnaD8Sxyrn5LpL3/+lpqzMPhcdWbGiWNKLkd1Vizk5frdK
/SW7+d4hA4Mv5KR7qcG/atB52OwTLhyvmxunwAGhlI/Mqd8JbyBYnZVPA9xk7yeiMqCfWh0pXrT0
EI+0MsOqCnU0kWOmmckktRzeZ25sE20gNa9U/SM1JxGeifDnoDjQRhhPktytMIMeX3fPnFSGev8i
P0h4NQz/ve11DfXrMNqxjYW6rmibUo5ogsyvl/QnPz/KINs4uzzJBgeOQl9aaUqpfUlVIM7UHcs+
lG+VfaKFCUGP3aUmTNtJ5hJt9UOlYoBCL28uFgvm/zaZSEzuyhB0J0WbfMwHqgO9taly97jnYbia
U+rCoxZT2w4H2cISnQxPrwSL6e7ONDC2kU1i8pIog1+cY6B3HuWn+/48JDN7jFGOZappJS2bdE9D
sGoe5EKecqlATNgXtUnssM+HqVB2dvLuITtTkKx25NTSl+0urfAY6F33pyJhW/lRaGPT8Nm10ivb
2xR0Rjb2x37/I/VSuqfTekzDv1tWHhN8M8W41copCKAp8AalAkE6tcm7vCxw1Sou9DkCmLjRCX2j
aVhgojWTShoK+zPHIaE8ql5XHEeoZMWkgE0XEqtCKaYl1OIsuqw/gBJmJOYWHYi6BhF5FO5Cm+1a
+MAYy6cKTFrII/YGE+IboMoO9c1XYqB0cY8MVM9Zn/TDTUh8JibtWjm014xFHdRSuNmxGJe70C5a
N9Sz4q7teGIeI4kp0DK9e08pewhMZNvrij4DqONTP/P4klBpvE04ZrJmuTE2zwvN/mh3o9O8hSx2
wPypTWvXC8PkZlXx3B2sNWqyR1MHd7VdKA2Dy3CPyBxzvQkaLJQzKxJStXxVSuoEeZ9vkKi3U3DC
NAojq1Rog/kJ945StEFB/flt2HwAdGOS+E6Etnqoud+3KAfWuUCjuROyDbmDAZXvVglK0nOBJlVv
W26IZHEc/Jmq4lFJVt+cUBulCTRyPQ3XPCNJBIFj4GQkYEZ7BhbDo7Z3tDorRO+nWV3du1ETqg5m
XH8h7aBdJ6t3A7dv/U1sBa+syNiCiAVGLMgbXT7m3N2Rh9DvvgVRQVfwDCUQCzrKYOhRgghAXq5I
K/JWtFxaTeSHF1TSdzLIcFPwgDUf3dL62NKXxKzmqLxG3sgiUjhJyfWW1kgQK3UlR2FDMEJ2Crr7
F03gbOGa9QCc/2KBwSpylOBhpWzLMobNtRkTjiu5VTfMfhugQxdKnSzUxFgXuqvdr8EEaDXhOQh0
vPzIgXn0eMi1kQdPYhZCP89hMB7hiCOo1JfjV3IReelt5TylZcvTfEMOoNWPiNUzLfhgu/W6/Egy
XK4ZpocejajUS7MV4do4v55ZiKweGaoG4CcvWLskxLrSr70o3jm00AirKlpP4LmqJxz5IbtM7na2
mRy4Vv1pHMj0WBwgU9hhPZXlRbzNY01oGwEKkyjsnua+0hGUaXG7J9kJzPwQxTHlQqd0PnHZfZMx
DkGn1Nie67SnhHJaNNIlalZTCemmOJ7pGQq8lu/cECxyfKMkoJkFZ59DQVRWXg+E5dnveYHPZiIA
1wdXn3P96LynDsIhR/+K+YvtxWl1DnL2N09Q5SJfoBuDHb8bP8aE12CpixSFRGg9lXbIxP9WFfz4
5U9uw7LKwWAvZ4yqMGjjtd+W1Q1fwb0OAPPhQ/pabPqzVY/JjaHeWVNVrgHIejH3X4J2/DfKwct+
wH/b3B1Ta1pQhIO8mao4P/+jgImnjccxl7iFkrW5TeM1OXYvVQbtJ4Ki4Er9j0BR0dOIDF15qVrL
yaTumD6lDF7h62We+kZD/JY9S3VlsfZVCCAVx4SZ4zDolJVk/+m99Si7u4XFlBGv/hpGiJ5U3ur7
NFqO6+WbVIbf2YX4CnL89nP+5dqN6LMH8lKs3jtYYGqWvnqvc1FSlujqCF1VvjHz3b4DYzylvg32
IpqsN7jliay5qCzEIHtYXOWXYqTM5/PwWE94hxw/B7WMs/GMwEyfTsv1XfMn+4f02coED0gRIjRm
XSIf/mNsN5uI/Nv0NdNh8ikO75fZYk6TrlzGuooLHzPHxchrcLY5vYhEgGPtbRYUs8D92ZBJjyNf
Y/YsZPdKd2Yzh/UM5mpJrSPWDRpxbsFOb3r/cWveIPfvuZozSbrJF1pv3V1qdOPGDj8JxywwYMpe
yXq8vO9klUhmTyhBJLgMqT/eq+j6t2M6e4zaz1uoSgF2SQCK9LS0rOuIq/nkr3xflkVfPdF9/pWK
t7+3xL+vN4PjkvO9v5Tc2TfaIplo8j0pIrLd4EAc5h3yC3jqbU9sewrJGdcSYIoxg2q5IQ2GLOxA
u046Y0tEVzocpotZOjVqbJY01nOKE5jr6oKMf4TlppGNhzZPYCgijRlglQMfMc77I7+3cCtZeSG6
odMfc7ajuEbm9TPKEI3X95pkbX/qy8BikocSFgdk7pvbH2JDrhJj8CrQZg63OyVrUctOEhE18IrF
iCNG80Wl0X8JO3P4gsilfA/em3c1EzaLTTtzGAMR8AYoszhU7GDMs8rZya/Vk1tEvHlNJzMxJC38
VztVhGm/MakyXelCiq+F5mifwYrd6pQ2y3F81zygSYJDF2Fx6GgYjyJR6b5TXYVN+gyg5LqU220M
aiE1qY/C1Rr0ErmlyPz0x3lsuCZ/MDDxgYPMhT4o1XDJvVrq7pzDm/Bf47GVHvPomHu41gJv4E0q
ZAhZ5s6osaC4c9Ldj/wPl+uJNB4rrzldMNOovsOAkdP6HOJIGBro+vWjoYaFAEaABt1r4nAUDE9d
VoP6XibF4d0woP0DCrsps5c7gA4Jot5I17i0BxR7tJeL5QjvtmfMGAVxz1IOjCBjKNCuahsdINAe
vsFD+OWOe6NxeFVHWPjy+aWeAxRd62i0J4uYb8NakjXPv8DFZUrcbIkqtvNFTUsplVTcK646Yjnb
2XKFiEWQqYmhMTrVPDlbHXCgp7EDWNsMVKigifu+Fgg5Wh8JOb1W0SpB83PG/thIHJypBmz2AxF/
23RAosOXaeonhn20mrLkKaO5Cc6IUmbGdOTvdRTNtSpsHVURFXET8xcpkWsWmRmaHaKc5gPBh7qy
AuCavMBYFWi3d/t4vNS0yy8rDi5fp3S0yQvDkdKvds98vfu5VkFOA+ruZyb7Y/nuMRfhEFdCuBzo
YY4HWp/i9qVOWg2AEF2XSrY/bSVXR4PE9mhb/q4Koq51ndvnTrSvgxHnqmxWXAqZ+czUHbqhYtM0
aBjyw+/Ii7fIsc6Y4hXzwbr9zJ1bJ11YqDWIazls37QGqvAIXmnjTdjSzHH6JQE3AdAjHBepIh6O
Y+zrw8E8MOteBBw1bYJjOrwQcVSzlXS+jSNGV5IFyPJ81nu5Fm8HkC+LAVSSP+iuUJY9ksGSFWeq
tLzgJV4GN4m0f3M654joomfPhnHbhUTSv2FZXC5mzLR66PMkMwdx5FHf/E+IceJOG0Hc5ln8rg9j
05eSpwPXPzXsxnMrntk1OPHoKNMtBlxjkK79eeM7soo5DuEMzTIa1wPyhVyN0tbbOTU57UmTTnkU
nDVTQPWaHgXJBPDyZ/XGli4TV5+Y1xvWxUhr4fYkb0U/a+xULd5skz7SciBPOvY5U+WWGSxt6vi7
K5CSbdljaT43Q+ihOjYfTVQsCigZq8v9vVNn2jAckvCD41IVNLEDBfCSEgzlGlD6kI9yjB09AxQ7
ks1d5UdZ0h8Xd+M3X+HOQiGxKhNVXAyTAYMacPUh9CNTZdOWm1+usq8XQ5rwHrvChl18nnA5B1qH
evTjphhUOiWa4Kze9rPsvfs6SKOjaRfr/FJMMkPkcJgxza4W3ltMYG9rJb0dMWYd/vqd1n36QF6x
wzP3cyyhSHHA/xyUy9DzA1hpLmlGjIG2l66hVGRb3ejm4GMi+BPPpZ/GSnzef5GDv9M60fDOMdBn
AFn50/21wLYW8+NsUhtHOLjuDsIeX0xX53PYUiZqpNldL0BjRcD/ccDKdvJK2OpQttX62l+PEQ2s
xlL3dsfgcNbWxpjjHIokaTN6v0dNyQjT0h7AiGmMSUQVbtuLlA9GxKRQLsgxuXrJkj12Yn5vPrx+
+OPl2SbvGQthg66lK/OhH4c/DgI8PLCnwpbm8pbM3eXP/PSAjxcjAd8IhXsAk0/pa++dMOeOoA+v
Z6ZASnNd4k/Pb89uSRTm7LlMjzLP+WFff+nLmspCxqtp0NXZaEE0U8tKp4EXwDduFd5VbGYvCBRm
gOPUWaCfX12MmfspDszZNnVEE0T7r6/Bt13Z/ze0Vtdu12nms3aw1YnQ1ti3vL5SWVwXF6zlh77O
Jx6DuF90yYOivz+DPczuHKZueisLpIg8W11q7aDsSZyoH0PTT7UtfVs33j0mHkDwZGdnd1yvRYhv
Rn/WXX+bpaTkbj8aFYat+sgljZxMQMfw2+I1yJyaMhHl5E6bqRb7n+vP9bkZUfHN8+VKkLRTR6Az
RLQHTvWKGalPPcIr8tMYJXRaw+X4lJyVnZned/pDevjg+0wCU9Mf3qphC1y8aZpjeqPvnlnpBQLJ
JmHTTGgVpiPh85Ff4InndTdhkE/ul0zsCo1OBc81RpDmRPWTDKuwVEKGh0omHVPYTVO/KUm2yRWH
Y17p3yqndNg21hMkZlh7Qlzt51TPtB4MGUtjv/EOnO3ZFrg0t887qS6cTfJzzZ4bOPAsPOKJngiZ
7Co64EWeSAui/wwI0+ALO6040+2B+YWSnJ1ww/pmxGWByPwrKmkuGpV6asjDBQHGcLZ8Eqmd+Hms
6V9L0TxAOSCUAq8xPsZ4od23kxERvIF8VFqXgYXyofNnVuyxcHqAGi/01SDgeXFzGxTI4cog2NW/
VAj+ZCg29jESAfQGavAM18hoN6I77/hc+l97UtDpXdLu33Dm73XtDvFprcDvH0RF55PlH9plv8qo
qG0aCayg9poZNPF7+SJkYPs34sqF4jbEQdGE/cwX4bwq7gVAZ+nt1hpb1DZ7wW0q1359T3SMdQvA
9YqD3S3m0FJudJVU741BFSSs1nOWI+W88+KVZ07o6JunqDIe4kgvE1HMJ17VMiSS1I6WoS587A8k
ZerVRRQyg9yDUtZd06lKuzkRHxmD7/bYmaCsFmuxVQbGgFkWIV+81xxt3p0MyS9ckWAceQ2gjTE5
ON7hXgBFARNMsASU109DMGiBVaWPHR1IKKwZjIWsl7aRdkWvwrkSAN/cRu52SauLoY9BzRfWg5wM
Uqt6ur4dGxjjIxXX5kD7L1aoOTMN2VF5Md8buchncWctjehsEtkDIvvbaDHM1Fcp4aNkxez2L6Ud
lBXbPfWLRzvgUkSPwmx9NtszXj4tyyTXxqX3/erzRCGmFRJ4546m9J/Bb2CGc6dbvgawexLTIax5
5EqV6d8gBYFkWBaU/sC0d8VyNmufR5xYZv6WroN9jwrrd60w7WZRV0rICQB/YgiJyw3ohKzkRmqd
xtOJEz8kGScoqFn72DhaoF/aqwMAGwD/kDNQb3V9CcIvkVxLqVfJSNY2VrcVBs29W7wU4pHyIAfE
vzFbB6k88TCfKnQq+q0rqjq6uShkQWzbmjQlWV4E4BZAYFxmNvfxN4AHL4VOig/fwbMdZxt0SYYM
X8h6D+XWXtFgt3v4lqecP4/0Z/uprP45pL7/t8byBhYXmY18N1Tp2Bp0tkk0nkJd81vMMgOS6QBb
rsTZh1+bQl7x4KK9buxap4OlBvuWg7uMd+6jis3gRaHqcczwEhl+RucgsV4BwbsN3e8kogdOkfMI
LsF1eeIqsOTxD5Z65Lv+IuAKaePYXVKcyM6s3bKFzjljV0w3yDaOCY56Npig+gXkgozGdnGUGtMj
eoGNd4f2iZu0YhQfLnbFl8mUawAWF9edoHQ58qAPlf1ks8iPiYgjN/dUicKOdqBp+QOnx6cLGFcB
F/vbcMWKsk9biYLIi8lRFkF6iODJZBZ+fYkwZUZ3Fq8kU0Kt7451WTpOYRl79+BhxSs8Tz9EVJ4e
ZOCRh/5lJV3NcTeaD84LXuOgmV5nf/qjAezPvUdhmsj2zte5Vpibxh2E+z+XNXftlbsviNdclMo7
4a/7teqK2KGiGOKIgpIRUpuVKs0k48sg2RlIS/dTqOTf46g2G0UMJoUHS6XwRFvQfS/gMlp4stFm
Wa/3zN8bD/aielwGfZFYT+a+0BhcPC69LeVhPzdG/Zg6TPLDhqJVz+TSJCAyaTrl2ATqvURQyQfo
Jr51yTFe3HZT6bP/ciR0l+Y7rPynfMXeE/WFcYsYScrz6IXHzxiRIeO4VUA0b1b3DZiT989y9sVa
LQ5hpfwnGW7Njx13u8I8t2tXho49CdV9dowAN4Ej5ACAdXG9Pu+1LK2YCdGxHYegOXBuPIbp/LEQ
UaARvAhPndW3eOPdvMX8spk9mDkK3lHO36oT6GH8nd/Jb+2HpIG19eypyNU1bIh08psUx8lhasYq
x7a49VAtX1/F3ATvReZjw+Ec58ExF/lli90KAcMcwwUK8vjT7Rp/Ic3N6y5nroADCgKL3ruhZfHR
NbmAv5G/7nnFHaz+QVBtpqui7oTjgAJqCTF6AdNU2hGKJq7wU3OX0A2R0dXH+rhWFnsK1WscdKLZ
n8XQUUJeUptmfDSwqJ2BUIx32/9d64rfCC0qdOIMdvQVTiUo2XoTRtI81lqfuUvJRr04RV1g017O
sTeS9iGUA7eqEXv1UBuURy6p86xUNHiNSLOIeQmBRzQj4mYPWKrwFGC+iHUmaIOrLqjSHGMs4QqX
mBmSO0NU6PuMCmyNLscVRACsR0AlQeWZvcmmf30nPw5NGXvxSIpfQuNKvEJlGJGlmhFPXM+kpPRS
z13NjxyAyf8XfmDsq99vs6NIqWld8gxkwBVkfY+cLY5vkbED+8PDR/VJZIY9yH4FyCwdnG5hEvBc
3dN5sJD2bUoWAmSylRh23t5/cCNpBACKGgGrysyD/TYTISBgiE+SPfIZ2A9jrolruoz3yN1bBypz
bdY9YfpkdkQBOVRtvJY7ZYZjG0lVegAFoG2y3str7famBrq2yUhAxeoGEUX6sZtDuK5zRGr8ZDDP
bOIOSrjeneT4D+nahUpMGVQU25OV+CW4u8cBAPCpQQzXB91bON7Zc7AtrZVtHvC5g6zptIZPXhy/
/p/6XjqmNv+EZdcZMvE87PabA7kGFbJ9uyUbl1srVv6lDDWWtucNwAyoWq7GTWYOwfjUd915DZxa
gDw9zg8Q2+c4pdKtluEQAoA7GA+Lu1D+p/S2nywAmgnTP9Tq7j3uqtzUFfJ3gpFm6kYCnd296UKA
rH0SNEinFgol+HeLnFy7t+UUaLLKYVHVunqC4BpEtJ9Myf1YuGGp8lJvS6x3w+4gLWIL5Z2GRcOd
jRi/ViykcXetPcGVuvjoweZkqozyKpXEL0vWILZoNRH3bEcNHdYczQ39mlXeEOdOWav5lJdnHMz6
qouX5S9C87114/jwxxiR9CkP3zLFxecSFJzQ2gdxb3qwTr/cvrFrH3VDxdeUH9/ZxjONs9OGmfjE
WufiNku/Gy9V+H8kPat/AbmAwWJTxK8F7j7rVlLqC6KpYaxKhRTm10nGzCV2/LcD8XT7wyrfZhOA
NAskecLJuwYS0i+M1cXy9IknCMsxVaVek3lmbswFAx15dMAQukxbHbE+7FrC2F6rOtH/4kBZ4evb
egp46VyNc2WWp+qLfEH75an3inkrbbiMYJ+yk1vKMo9grY6ghkrGYrpfTacI9+vSb5IdbBt3iG6x
F/KLLmdP8lh7mpCkwyrfYN7SfNvIprJPW9eMCRVqX5gxTD7/9MPH9VQYszmSMWRsqjaXJSkV2Sqv
iuG/1PeuTfuLtnvNgVYB0vbeu7NwUh0cZGjpy8bea7lcCnEgj5m9Zz/SLNrvtmyDRkH8yKCJYMkc
y3pstQGPJbingDPdVoWDB/8t3fHNw1YjdGI6cTog+TJgstee9+/18pH+8Mr8qxz1nWM0L5R0vlB+
4zwsS5CaKyERfUIGAFK/wfW7JUm/AB5D1m7A6k5mpNdRd0LAUpP2Tzyod8YVuQ9Kj68Xst8yQOYn
GC+c9CfbRucUyPXPE9k/FNyX9Bx6AApVfWYHPYqRahZ5/h8F6K2L7EUJMBvosXWtfMBAZY86jak/
BHFImEGmz37RoZBp1Ydz2P/MraWsoEgPytY/BpXHSvTdT0DbuJZIE0TZghxmc20K4FziFBUykb6G
hI2juculU5RTzNZNi7PjUtDSYaNn4JM9dn9k/jaTAh5tiLFM58yZUmqab2b4Wp1wPOXiqCVPGPf3
GWCb/DRl5ood4167hQ1djpN0/u5VXmb324+Vs0tXWvUxfJw83ScfHwKUKXvS2lMaQE4lT3mu6KCO
KTKrEeqk+Ok4K8eHO4f82JAGrENogwzUV1jx9E8VfNhf28lhWQjQ5W1/A8jsPXbPBJ/pu0VxGhG2
zcfeBrPXHxIdovj3m8Bz2C6Gyi7OcVslPw6Z5+vLgjmlcopCLVgO1J8MF9Bv7lTePLy20inqe6vG
TxOM/kwC3/bkj7SIQVVx9nV5HA9sc+ameHe5NuomDASSIVsB54ujHJi3IA2bcRXjI8zh9E9Ck95s
tXd3pesN5PUxH01kScMs8o1oofQHCJQ6bXClsD4YZZpDEj6zh727+FN7ddSg3aFHPh2an2yXu72/
1WwDSN8pzly/9LEYNemggeRPQbrKwyj+sekRYod6BbsB71jaagwdy8ivoNBFXyQorphB9KGdVvL6
XkHDnsIFdNBF3bKTwAhBuFr+QH9Dyzbx+iBb5bBHgWsSrBT8xPVsM8uCyW1IqLPo2tZxsCRjfvpb
xAdXg1v9b2dGspmcqlhxuzG6LXKhhCf3sC3I9o2dZBikTVVt7ZHJRiqwjbzSIa2J8EO9hfdFGeJ/
ujzc8ZsyyoOrCohXIQxsPZLzb+wCyxpALoIHcJnXI9Rh/DEHk5hCLENhYMzAxLk9YjCGRUT5zqb2
BHQI690aP0Q0hLlmL09tNaI0MWMY69b6WovlepSpWgvsrknsZJ63vrFxGXhudNcmXwmOw9lLaYE9
boq4V2GfuAWSYRqd2Xl5GJWjr2uWrXbcj6KHjYMk0RHUYvDuyqqBeV2S1lzZq61a6Eipw1rJTMv8
sXyMVdvu2Gq3oAl634ykGRJx5FtKOjYo01JbNBYNGR3Qn4kh/TexR8UUirD26icKLC08BvWnRFMN
xYzi4J36L2VHLWesjr45RF5g4zZz3kdFlivHK7hDwKDAPmJafDHeFoq46hS747g/sv7EQe5xP5v3
EkWAu3P5vp9q1w7crCVz6VeUj0Rxilv9AjmA5OgcpT1E1WV0MGMqcAadfQPzUBoMyL88MYdQ8n30
LTpLzTwKTtKEuCN3pePboGuu3Q0+MNRapXis8S4dQNFO2bB8k7PXth2Jwl9/Dyu7smS673bF7Dow
t1fQlufDXAc4ILhk4EPnobJEl14X9pDyDTDSLqTrv53L2JAspMlIQjTcEAPA+teH01tzZHWaVbVB
B3zto/ZDwhLPEKFTGPbIfQMQRY8+5paWV00sL/mooLRdtQivXj6Ro/tV7iBx9MA73X1Qf+ONlvlb
THLKOzkyjRLzwQMXC1QzTa1LYn7Z3oEa87Z43xwXMOyXfUmgnTTnsFR0ESjaE2x6KMqbN25sh/Ie
5Hna7gT8i4QempAfGwFA+GzErhV1oi5ZU3fnEoT89dqQJkVsgsf31ViZb9evQu+wEo0EDNiRdjnO
hGoOJFSweMIURasJaNjmzkktdEo7YmkMvAGBLJyssT6IV+OiFRMZZE8U0GiK9sQ65jtz1Za6YEEw
mRNZ/X15ptyVKqgSrzLQJSiefwY2fRNuB7A8e8b+rrWgO01MuepMIc2Nwk0iPGYXdjHAVzcD+Uzr
KAcyqJjX3WYms/L5GhanrMYUQlklYHldn2yQh9DnNzdII6bpsMNWzRGS/vekK20FCePTQATjT43Y
bHTQsm0R0Wp9FB1J3ze8zuXuaQfaezLyI9ZfwmwQtykA02T8wbc11aCMnJwy+K/6DJeKLBz6oO/2
9q/lZ2cdH6HWHPMXqdb0TsrSip90sFiAcdyHw1pCVQ7OttMJ8HPtw3EGkBsuRhv/Je9DUxDfgxn7
ubVhU7DPWdyV9ETjtToojFfdWpfd5AQfWtf8h6EiOfVVXhNzmjjuA3aYv29zV2zLJMomVz76v/h+
JE0dukSuZJcbU6uY1RjLMWV836tHdsriwXXdI2OLioSVgkSQTD8rMSW0SbQPEqJsrwgDE+wcj1Qn
GLG1yzOt9COyJVBu78NnHeGj6FXJvcYlbEtbSX4bkAcA5fR4bZoKoXJhTjb5d4Z2ddPcS6/Mial5
217fGPu6YyOM+CSYhhD+BesNpUwnx1QCG41Q7Z6qhsisLWBxbh8aNb7m59onEj1y02h2IPPvgJwS
pbVAeKOb2USj1pJcoc6BHeYNdg9cRdhJLjdL1GPv08KcgCbUCzmJG3zNmkdOXAy45q3tK0JaQ6gE
lk5WfvFCeXOOH6yVHsp88vAe5tfk33acjL6hFRtFdw+46sH+/I6q59clGgDykWKUMVRdZY6ckPn7
78REMkIk5xVqNgHmfR2mUgGL1H1mecrFc3bMlyIAmsB3ca1Q9YWCJGraMfvEjHlxTMd9jDtlilsi
p21Fxp440VvZlw2dNFDmoegy9zIDdJUZ+bcnY4wzKJfVqrJ7yJ7m5xs/7zkcoeJEuVpy3+1t1/Fz
7g+fCIFtLFNVSt/3y4XMxmZn3Dt0ildSH8eqDpBbni6162ySLCoIzTqEK/zbxcTtgmTIIztnhtNK
vGKZffieOaOUcR80Og2UaqwLiNGs03XGYcb9Oqb3JKi1qc3gSscumsCtj5nmtnivzbDtwuaS3V+2
TEGtd7MF7lhgfvJ2dS71i7KyREcWUB+cdeeR2WSzOJFa/R15WP3v97cPkaNhC0JWvXvRZL6tTDdr
Oh62iCkPE3FJqiXdhwYK7KHm3xPDoT9NMMw01WY0G2XVSWS/iCaiN8pous8lcCmtD79mneFFl+wN
jvxoFsig+QJ9SE2k2PpmYVNHxGJTDWE4doPPRbe9Eohawy1d+k4fsoOAyabt8IgPROzKCJV5URUr
+UrqCcmnCZBl+6/YEcbhLOaOQzhpSRv1w06DMvTeaeJHCEG8mgKxDPPJf8ARiyhiFzrgied/oUly
xFaGZl4q9wxL57v4DWgcBf0nHEl9RDy3QY5fIE5RkTJguTXgSUVo8ZP90laoXIbGFv0ZqgHBeW9P
TGN3rvyxec4QRPipMD54SZzgLupN7NS1K/YsPEI+K4XrIcCWNg2jDCQYBXaXVDEgaC3giJZdGwx4
Hdl5qHZLqy2NVfc00BZoAAWQq09u/WTYWo4PCyheA6MAC+ha8fmoV8e42eBP8H4ZxldSx8avY1BD
h/4uBZvUh5a2Reeu0EIRytyB5YT1m6CRVOa+iXRIonFYmk2Bt5Bhuhw2DGmdTjl6LYIH3eua40gR
3FoRBJVh8wDKUODApKW/VCAmWWFXX0yxGD/I5uRwHQ4z/jb5TXk8EFcKpgcTxobjUjzSW5MQmaQ3
POB7ect9XFnH5W6wnW2tgD5SFHcgPNhpsilNTWpqAIZI0Zn78yhG29AxVTveBu2pAOx0tIvIkPLU
dGRN4ovWoKfmRa+KgotTZG9cY941BKtLbRUfxOvabSv71OFKHRlsj8T8qrmVN6KdjF4KTXvc6+Ty
fysBguBilbN34U1f14yLEFT3N4JsZf2avaIV2JfJuBqqY/HilbYk0itWNYvZXpFQe4DceZBtNXK3
XPn6dFhoDX7leEK1kmvZdBjvnuj+Sbq54MDwH7wGYLphgDTVX7fbnpJk7hK+92fYjj3z67khZUGu
HLNF47oUSvYeXogk3yJWImxwFExxFfUOJCaCesPQr3Qpy1BxFZnKKa62g9wgn5pafZDHx7VlutBb
wec9rngZs9KhUvlVgsMuq06CZAZrd/tA9yRCWFQc/9VXAqCYVGIA0tazhy/W74Q54pJkrz2+LV2R
vWAsvv7aqEZqYHafhVY3rcVqdjwcDF1+Krt9OkTvOhL1q0qJSIG4Ls9aLmxRfZJTfx1r9fzEEzKX
cAHnuIx8rmGaACZVondEqjnS24YwGEpDQiMZ8Wy3aXhAtrCCvVw4ry6/XNdzDEvrEcH/Z96L+/vE
ImWUrPvd8q/JoxFWcizAZesKgh5EntrIvs+lqwGlxyeeWQ+1R8kT8fq9zLiFm3F+mg6k37A5RlwT
ZQfbdUCBU5FEk56gg/X1PKOf9A3J6W76XgkrTTQGTAKBabfZPQLAMdqAXPAF8r46eerzYqgqST6D
hUaZihmxhlhxtWasRCt/C6pbZXspkUBRbuQ2yZkpn7B6xke27K00N03Roiq56A+BypD9PQeGD/O3
0dPK7dvYJb429COlN4cvB+IOMqdq9edwLdWEF65/7VT5mOIbskTNbbpivZcoaYjxYOA4Al49/BlI
lnxZK9qc2y1ufDE5g5BUvbFjCaMFCiw9wsljRYHUci9MK5CPhXCtm+Ck5OEgk0kDR/27tGeDytot
mxPNpRElhIlJTb6jYR6Ynql65G9TSHh+fvLZuxYfmCx87cPI50EfMdF4X6/T6Xy7FLVVhIZsm+QI
WohcpQ8ejmIYlRPnS5rVnfOIQNV7iv+6VlhcMD6t2/LOMnNvvdkkfxYv2/n+SLVhfKE0FDdN1u9+
9HDPgquaziRdLpEo+I8qyVHkwZ68e1g7+i46iZRSqik0nB/w4SP+Z2Ar+OzGayETe0IACSMWdVMq
Exr7lzCHID7Dmlhc54diz3GhJSIuHtFGwb68Bz3o7hsa2VZHGs2RJjXjQLj1pqk/v3qX3tNwWrxi
ap1bxoBIPohfU8p18xBf74E6l4TJQG74jbNm1jF2BlJwNj8RoI2ZD1xjcRWhMXT8XvKYP3a9oWfS
p8H64ELrTUuRrS9NT3471hEzcUw6pFdsL9tq8F1eaWFPS0YylhraFQlXj9t304kLaTPb7EYvGMDA
PSsFsl7j4GMFqMPYLJuSuZ9NlamZszB/uoDoZoL1BifQazOBcw0PnuVb+8KDZbSaTgWl+2g9Ky6w
PerNZPT0BF5iIN2O/BhlJKpYcDhGDtiNipy61lXdizvTy3ssAa0KQo+nYHpN+71yT/yp40rtezsN
XrUFBBaiqqKoWQpxvKV5ql7OWp8aLkvi+hOnU3zUWOFZyZ8d39lGescvHi3HxB5H4oT5ivicBRZI
nTnR9EJp7aZgtfOT7vdXtMOfU0yCQNmfFN0kbrrkmV7gz+gOydsyaDcp/IXUNJV/CRAsjnFF6hfB
l+7U0VLCOpxy9WCD44pMLVdc4tI96u2qd4df/pFSGCqflw6ZxmIUR6mbE4vEFBIukkNvjcXaa5dS
8m2e+z6pMomqeHPwS1mjW5y6nPQEzwsFa+5W74A/+0WbJ87W5zx7ESeT6g5UgZQfLptugWH5WxuQ
Qc2xGbFeg1tVrjZ+pby/Mo0HwyJDg0OyjEljPPxRD7eODGb2eRWMikY8DkBqkxrFlleyUsJ4uR8L
H37YutxSuwczKpRDQ+ieFJW6HhMa/jBlPfy5cjdLMPf27hVi3WoEDx1AukwQ5lOukPcVfdZ+gPs4
frjRuD0ho97zNApRZrjB1c0q/FpUb9gnNMo99RfFzTyuCn59XF4wMkswjMbwz7bZK78OVd9OGxPU
SaEtdaytoMqMJuX80E9lCpE7+jO9J62SEbzy0Zwl1UblBVqI1O/pCYvMSLr8v/nPcbSeYAr+Zrb2
Jfs7lRatW1SVH1ISQoWqEs09Qvpu2WXcPZG5sVs9jyYPvCDUHAMevnOgeByOTO+G93b8RXVlU2Hi
XDlmNe2Re16QCNn46g1XzaoBeuM4v6uLceE1UxwH6+ZkKQD+zTVj/YRFXzG9TL5Ap00E283Y0u3n
NpbNhQt2w95isMHCS1aDBN4R5eRqoxgK/0A18Jqisdu5CBbAEK8kWwk6TdGUkm6IT8/8SdYqCX3F
S6o14q4wfuN9wK8nVnRv0ADCgVEe2G54xuyyiX93nnP/hQZWu6+fj8azBRcjdM8hDWik8TMOBtjy
haV2weN1xCQ5XQNCUaaXbblC1KOHs96P29ZJMuNXVTNcgHpWvd4I02eCIoVNYDzj2x/vxkD8cpJu
m6YYo62bVf5F/B9sYPs8FcGOz2qgz+7UBkr5UmtjHnPxC5fM3qIViJWjAFZxbKT6y2+7/zsr3ejI
QLPKcs/s0TqEYq8Ri7ydHL8Sxw0xRLfxnw3HLuYuAEk67EKW3t9ELQRSbauCoedJu5o1LVaT3neo
ELvtyH40LBWgYzXaRDwICmREEncZweFFwcBGKSdMGfYiHNL9zBNfeEsEbsy9nNSV5v/PNfy6B3I5
5ZOESi1eJGNdpVQHGBAhHowPD0Wfg/g/GtXw0/x9LD+SmdfcEu5P32zxdHv3intnJl9wi06RQSaI
geLSMoOhNvuXURbpnTJHsObBLimDNEGiw0byDu22QJZtshjg9QY5ES68G9suITPFwAHu4zpIkJGU
MgDH4pgjRbOu6RgM9xZXuYjPjLHjDaXKAEu3U5lMBKbZc9TF3OKTgmTY3FPC5+p5BtYOmAEtCFuj
ynge7FU07GL/W0jCiuWAiUbF4Blb0xAt9LMnx2eshl8RS7v2GgPPI4r6CYrEOrNJ+cV9sz3284Wt
X3UgQG3+rPU7fDA05ac0+5z+50qup96cg06YEUlNMVuMzkQ/oporEzxk1htBazSBzmhTOiywYcWG
QzF6PLjAYq3YxiSy4vZlgjGKjKZVuOeu0ACV+TFuIm2Bv1xFlSO58xnL9I+jHRvARx063/IyiFTZ
7goG3GWZjsIbNkAErOGIS7dAzSUiMjV6tJzGqI+QtDyJy0h2fsYQvxy56xp9d5Wqovlsdr4wMzHO
wpQuvPGHK+B/zG0JvFTCpWHhG8l+FDYcR+up7Rw40tZWoZZP8reY/QLnGS7Xm7f0YJ94AFqrthLJ
IEjmVFr0B4kyMpZidG5/ffesRkV9ZcS6qFNRSvSneHrx0xBTXdnzJjmRJFGb9k+bsMiV13H6UFh+
dqEVxHLmV7AlXncwksxAHVN8U2+99wFXG1OGraiGt0CGVBo+m0s/Vmuo7S+TKERHigmCxoqRnETK
OB8jvMuKnWmtZL+GWXi6svpD8wwCGI0SQj1wQLEr3FfTSypiSlTuUgBNq2Mots0voP6AZfrixIYP
IMNRsbJSVw8qEyggP3DsOEsAJg1Fg0Wu2kQjgAHPbw7JC/TorzEo6CrxAVEal3/Y3leTcTYoTnb8
nCV3fcLGsirOyT+/q66uVe2HVy98EvRclz1DNsbr9ZRflN/mZFy1GTfBNhWTfpJ0mC1IbLvLF3d9
1iv1sqrd2Vb21vS2wF/qFOL3iu/Rc4oCdkzDNcv2inFUrRnQcHDg5CfmAIe8m4fp/0aKBPsCZtan
cM3JP/40cs81vGsInIRAh0ZaK0wGbpDrafB/vDD2Z4C//t+5MmUMck66TTycRwlbxFEEtt2urIFo
U+yWvVdS6Kw7BZiye0UTlammRJgDcGCb0t6FBgawmK+HXosDG2xuAxtXOeyL4GGQ3XIfQJvzsfAm
UMQwBSgvVh9NeF5miCAh/RUnwqK+KEnTG0OG/Hw64Gwufay12MZ0cD7+8jZ8/ISIqP98wD3tY93k
l8pWK0crB/fCinACaqyuQ71ieHuzKN6eDOzwBEwioNJy9C9uoM3PB9QZehRlOCsej/XCP9plBBeK
fbVUMnNirU1J4oHZo639pR7gWp2qAL93FBTEthSDQbOHDhURzqYlWt//uk3GAVWf2/PCfH4bM3Hv
du13YhUEJJaBZ7uKyzWeUg21YzG6HJYcI01U3pHRiu7eP1O/gm3w3O6E5t02kgED0VclDUM+kvQb
1M4DZdgzG+h3TL9vtv6rMpbwjkXecL0YpgyiLcwHLdNx/XJ+2p8eFJJZ+14LjhdkLmmjY9+/nepL
HNqszeDqFf6WluQ1uGVTdOwN3AFdH5x9uMFNzUIGnuIwobn67VUB2hRUkPyKQ7X2I63VYMAR7BQi
ybCLurpBCdkX+maHgU67hjipwZNUa0hCJcnIPN7OCyUnvAS8XhtDZz0xJlvAL8Rpn47Uiuhb7VhF
wq+0eEwCOMHmYxdYaN59ybwioP3IqhQIrLsBIU5pEfwCit4PvisH6wKcCbCgDDotcr+H88+Ge2Uu
24j76OOxJbWvbVasOHzrM0VKXay/ior5wXuYbVzTzlZ/cORG56TeLfuayYzWZCDDuCJq+nNrS15f
6Hc9B6fH0hJI1jy5QEkDvNoj1PLrF1XL/mBH/xX5hVBk+M/kFBQSoHDYoUWHkrjywRnamNysFt6D
C8ANfFfROyV2/ae2LLhaulGBuzaK+aF14bCX3bZgK9vvPDcZUX+PK1MmnwwB0OnsHOJP4VHhlBvg
Abq4/aA7EiYhLqwMspQ46mfodM4vWP8pDDtK6cltruhyf6efUUXtjmgCr7HY+p2A0buMtnsfUMyZ
/7GyvEB8k/6OUWKQNO5UB1kP/HhxIIUwZ+fuOZPjxJZLjdv/Cj09Q2m+J9M/EAZBY9kTM/P6ATgW
9plC8I+FTSMxNtIhju561wEn/MQ1lVxzi3uE6Pr9Vp7HfZypzo153x4ivXQMTBVZUmiUP1v0FTEA
mMDSUMMnnTwsrnD/SM4iUI1TE04/8wSWB3/06D8MTKYfTjL4bbZYc02t6AGE8qSE+KrHuwju7zA4
4vgYU4UgWDa7l1nJFoHaFqzSktF8hCCiEJru5usGt8rQtS9hjvzOzd7X+6ICPQcUzSom5ZQGE5Qu
Bb85vxlD6MHweKVUAKtYq+38SDeA+IKuQRgcU4/rhnjXY7LRAjaIlPVjwAh7MtUkFxsNSsguL/eD
CvftdkCd3eIFJ5FKFkhNl4oxiTmQ1FY+ih5L6LNZya2ZzlbYPVL6wVqiyVeWaZgRqDs0uVjgviAg
IYQUwEyJCIrN6UbVD1w34/xEKnc0Z044Q/tw94TEoeTF0gh241rwPaLu5rjdUy+5X6cn53wEEtKK
FOWCMcOJj3YLLrJaj8FfddmBDPI0Tz1j+R3cbExLf+KdmvrgA6UpwZH3xhSvnseotfGr1yKCwBeY
jhHBSeJd1A8/HrrVseayR6IST5laEJy2xpYM1bvY1f+XcBKNPlQIImXgVoc+0nz+AnvuUJ2Vd5oO
8mSc8YKKaSe5dkaNTU9ZWGRF6zMXnGcTvgiHBikG2PhrS+uAI0ENENHvClQJwkQVw9FwV4nb8KDq
P+783/fDu1xfGgqsVAHXJFwSPWOAIjh6cb6ZF8N/OlkWjVV9twQIXNfpeXuyCWToyYSnOsTt32+J
5TErbUSwXpJquLVjFyv5929uVwtKoPN96TYeRBoRvEv4FCSruHdWxUra8nRrb3bjthVXhqoxD9lZ
rsovXcBAK4XmVItypXDAnbp537j7sYXqHYYksa8Lq+Rd1iSMWwNfPnSo8C57qoi7KfkQfrWtuct5
oyHqw8B3iPdtkepXsfZersuoD/PAXTt4X2ED7fXJcvtod6thUz5zEw71HoUda8Lpwm8hMTQlnsu4
4JkCXMmPWIHDXwyu879JYPh9ENpKh1HSWt/oon43qEFUGHt6wXzztqw78ecqH/uREOTwUcOZJUev
lQIswYzGJjfGhXsUEVOvKjYui3y8kqr46nBPiFelhgdYHIQHpQcwxXJlg1bjXhkkNSH6aZn6ufBs
pLB11jM2a7YhLx3Ql4hSVP+sIAjj7qDMdZvlkdd1iIkNyNI+HF5U/0YCzI5n90YdavpTG3ZDJ/6x
Mx94oaw+h1Ip8k6V3Ylr32Gxmo0u5VQVS5itjN/6TML8wbzQi2KoZtuNJXu32erxCvSlFCXM9tu8
z3MD49DvCtyFgGnul7NXIuq05TDfuwpoZPyufMH43Uddaener39eqTcLPdMcHt9O6ADSb8+QuOAx
6ckjD5pEK7v860b0PXhq9KzhYrNWllbGpwZo+wM9hzXQNb0lt2llpVd4JnZdHIGJ/lRt6B2JXeUR
vutnGdFBmCVUE4W4e0PtHXNBup6nh8KEdM8m6g8/5RdPdgdKudjTsUadBP88gbfYzm6cUb7rMXI0
sP2Z2yDDTMscLRKT96BAYGa6uw+gR4Rkl2qQ5xSL7jbqQGWCkQSGuPX6/Z8qHCGswV4RnBWG0Zr7
oJ7/TDpTzKI+MjdqLTNajHLhaUwFCAfjw+vsydeoq/Xp3oveOfCeljQ5FHlEFI7EH5aUCsOl/D3w
DiATcn28bvKs+Hg/+3tq1cWV0IGVY6NrAFaY3BlhAP573jJhkFkRZmST8t2W1yI0zhLf8/gq9Lix
So5Z37oMh2eqPpBXxVl5/LhPNZrwOhHS7aTRhM0Ggm3xQR/UFYajOUgAO4f5+tpQvIZ9Sv2cVJ39
R0SWyNwMd7FW4NRPuMz3+ZwMqU9Dx3Z0QXRInX48vrTLaXQhCZcaZ4CVvBv8ppQJaoHFpbuTb1Ly
RL3L3OW7cvOVzChTTi3ap43ukWuXwOFeH7xi9jPxjaJRY5vHxWhJv/ZQ84DoBVZWy4f6fIQBkkvy
+0BOdovBUjs4HlI7PKFLgKO3UDRh79phpmH4Ptp/ZUw0IsX15SvA73KsZcnB0uThaj/OBFAZusCh
ETSyW6M4G2+uL9CDoHIx9nxF8e2v97E71dtEvf/tgL9B9F1mqCNqU00iWe/GWBcK44bKV4WnMIyr
mVA5BB/+lVkK8bLyZMQ1MLmtGYHcRy+EVSSFnEhfatg0PsdykNp6uUJLS8Ko53J8L5rq9ZhC+0rL
tFaN6a2OdzxJYyAZHrvIc9D4B1qEWWL9T0wQo5VkbOlKcK3lAVyc1OWlGsrCicCS+FSxKtP9rGpG
1D6MGkD69ulSUjjkQZ/4jLWvkGXb3fJorn7v3BLezQSgg9skoVflr/o5jKMSifmWGNHZ0KSRvEDV
yYsDeKwuJv9PhXUla6g1YMSG2FeINaflUVyVK30o6iJCJDUDKzqIucC4gxtwXqbjCDkgag8CXGY0
WjTSu4wNu4I24pq5oNsCM/Quf33t1sUV/csMw7hz/c0TbE72Ncm3olULcYrnl7MoVc8bYXDzIDY0
yYQVcYYe4Oxt2+Us4CU1L0wcd0kChBgHjzL+5NxGZF4XJOlifKA1vVBemusck3+wrCeCxdCj2GGq
dJqmwzES45wdRoKyWyN/S7QywS0Er//1A1Pn20J26lSuLcAxU0+ca5cC1fSwyfh4tREG5x5KvO0K
IPdjzU52rz6R27MHJIj7M5odkk9I/+PM7hlfbymMaemMe1J8G8G7sfLY9YtEjZ2k/UOulvok4Xrk
qGPxyL/cinJhmJOzWvHRr3CuWXT2evfWz71PtNTlMlmB+LQttVKP70eweZouPA2zhrBQLeQ+KOgC
vSI2G31HfHIbN4UjK4pMRLJD7LRBGIN7Ldg6f5mXaYM/rM6lxF4I2U1EVJ/014Z/esxTsIhPTtV5
OxpPxmliWbG+nVjGbgQvFnE6UPN/XMaiT+vdd99TCBJFtjmcVweFcej+rCReC6TzHkTJs27sRDEI
k4MZ10qo4hch7OApj9lmLMf71nO4xlOIKCh6BPRTZuBW9aDNgl1MOOBuvqlS5w8puZTotVcCGBNm
uTBdjceD0ZkSYC3A/ir4f1AByP3nA+8+yoxkcOmBY8YPD8/ZZdZI7zVTweQZACA+wXiKj3RMlSXk
qpsuDGI4ym9qmAEN53PKfJCoX1Vbvx5JnpfUIDUSZBGch0pIElCqUzGnMVWM/nc4FWOW5arqrlnY
G3vwFEAuydOR9DlXquh1S/7uCJvsoqhOj5laWNXw5LBIzcZ/NN2BdBKJMNYc1G7oG+bPJa+Pkl0i
6hVvHoVnZqwrxQWzZytN+MGQ1fpAaTn3xBNUuHEeeJzxruTxDUWvdY1LRolcFMn2Z+NDXANcK0MJ
0KhhUqKKtXiT9fUV+M26IPZIB3nvNRp1RHIL/qYW8+e1R06C96RQ1yXFZeNC1cHngGCifFiC+3RW
zQTNTBllEHCG3ygXwdV1A2zdKx61OL4bYZB9A5NzwNozi2m12yC+nHG25wHOLmNPFX/AoK50U6aP
YGnW7IDEe97AlKS4adZaVwZNSVBzTtFZ1ykq0Zbev5Y/hh5zQRl6wo5iluaPwQTjDLOAMN8/k6z1
+jpptmj5jA3MoPZVNa+p4mdX9vCa3cs3HPeO2RcforizFX4kPgNJXeUf+mt21OhZSmg4nRXoSC1o
bXSPnMIyzH7YEHgnrl38ZWdRwvdTNlVVh9Rn7VuZttFvniGB4ZjSDquw+NsiTzm/X+hxAM3/wOCW
wAuqmT+HjRL2n02VnUvxxQmxEnj2U2lqVGlDL7PZ62ZBoqdc/fAsQZqgCnvfTZCq7Q2gbcqqofxd
SUPe3m4zcohSTQy1keZGETZxDD830C7lZLC3yf5LKIlWKIKqj37Q+y2C/ueJdSwLWR/8iHc6697i
TheVwMR3NCvcCjmFrveIT+70EVR9vyK2r9sIHVS5X3NWHEhZwmKiLDIKoHLYJ8EE4K0DGCLU8DQf
/iyC2Khi0AMt1MULN5H3hD31buMf2tqoNXlp6exHDR9G0EL6kRzrx2Op8sEGz+mQbSR0oc8wSnOK
XuCRyDvhGPuAE167hKudR5ZkMpd8PI9bCJlmDxFSzldFIB0I6SpiuDNeD0QQf2vZzDZecnQAgGc2
PWXMiSUoQLydg/KEXnXPdW0Y9DSxREDsmePxcD3tNM8tvCo/N//ttUUIefpnqN6Cwvw4VXF+nhGl
82OEXVX/kGgYhiOJPMeBky+wq79pDbrg1VEfvaZbOHUg3r7o3LnVO+ppsz1+OkeNhFrcVmCjhfaI
yUMC8MIUAHiF4FVK0vviE4qq5cjiv0/o3EF/me6yGoJpbP2LYu9Y1fH5AiunHPBvLeNwJLit3NJ/
2ji7kMIFQKfzdH6tRLUDe0KNfVlVcpRuwSzBghaJ8iTZ6YsaNaFkCdPCn/sHWyq0cPvV/i7qr0sx
HOzFw7fL+5XV40Yfy88zTzCj1BdCDI6bP9pzJf6qAhvMz7T2WskwoJC6A168sKQCZ2LkBWfc3lcJ
tsuH2Ab/o20eXIEstUsp1QU44h2EAyxepjiGdZy6Z0FAbMaYk3Tw6yRlg0NLrh85E90RATj899M5
xLAuLyBfqwqr6E4pUZC1eo28SOw2dnkqltpsMLuwHWYs551objYOitGK04+TA4s+R0u9hsufBzVK
EukFc4LJCMZyK3CCkU9I3fz7ix0JoXj2aGmxbQN6PnvgE+8aQChowTzWturuEld55Oi8Rmt6QxFB
68SCt6p9TVITeVkNbi11bLFU6H4itF2Onv37G6t+BVMdoB96HTyNkeaW1+P0lgB4r4bri86iDFw1
iORt1TZxJt9RX0TmsMv9ehqWuZEv9Nx3sGaQWC/2pxo+HQ/SJK60Ry96XXzB8q22QqYIimHic4u3
8uE+UXzRS8/0Fm/MqcUWPFHI1+NPxL7LymTb0u4JawXpy6jUDW2Mo+Qf4Gjmdshua7erMVjAZBhf
uBY0HeFXV9XOwdDAOeGYoBQbxbmUBce4RshnzL3r097Ka62y+EZZ1j/jKREZsXCtEGwGicdgcyar
YCsPA30w4Z2xrimj8o71+xwGtEYt+lbGztB6ushJBYwKzeIpwmHdOraTq7I6UrRzi4/RhFBdr+d9
2v+gqLvXwQ3o4hyVp7g3qIIlv40z1BOnCbEyEBKQZXrtPAfa7PJFyT+cTafgWqTZmON4ZfGF3pU5
b50AzdC+Wjmi3NTdMOlIIUN8P0Mh7+9SQ26WlNWIxAC/1CpM/NUkVjtS3mhegURe1PNSYDokv4Il
6IStzu5VT2+l9g21suSh77Q6sA1NggTZPwvLqw6Yrw2WnPtx0mc7ZQ5gUizOeDWRfONmujWHDAUz
NVvi6E/f0fqWVCGsyrVmZRziv52HSYvrZrCM9CFLJ4oNHOVjeNiHhwxvSb3gp+pPkouMOjC/hZOW
LciDkoOQF7FTvmPGi9oa9yaBcmHMRpN8ijnU8s4BwBs9YBueJT5hhp4eAvvv8QgxUAYkIgSfSgrm
ud3fOF4ECD//u7vwM2jiCfwBpS3vmGztsjPnXy6pbGfoJF+Ms8gDAQXcqWjrELAXf9s3uKG1+iWg
LH6zZJk000+wQzoNu8TYo3WDPo/l9w6I99bOxi9xpzYAwvRxm72iuoG2g/0o6D1S17e3DKF4hMM4
Zi+rnXRbzK5if/KPMQcGagcXMQsvrPGrRg67zO/zbE0t2MVVZBvqlUR84Ulr/ApF4pb6PD/6Np5d
fyYoUR8kXhhGvGlI7X4eQiqnTt9od1cpgXruxTnSxJ/Sz6jlYAO3iDFzgCEwHXuFV5xxmSeYzd3P
86HbIMH3zxrHjETShjatHBVwQKfAceQhw7x5f+JkcVmWJgPPIKgXjs19MpTwF92jWdN/CHjvgwYt
FwbsmpUI1FU4zUIdGBuYlcFwhJF3J45MeTO6uoHihN8kv6FnMqenEcjeFzjAIjfd3u2fTmHwshsn
zXV4DKUyn9mGPxMlmLyX3j8lspCaW4EoE2+ZQnfrQOqsr4b/Zt24zTKT+ROaN9s1Fa/QQje/R7t2
bHy/Xn5pXWbJzysTvLb2Se7TKUQ3f5xowJprwu+SpqBkcC7+42tDOSBBMvrACCkUf9Zqchwxgmty
A5Tvn19FjOU2BZlZCJEdH0peOVzrfLmp4/leMZazirjbStEVPD0yUZwXFeo0gDIWNzHRzZdMWGA/
eV56kFU1uaj1hl6rGsS0foCNsfGbHQuggSjttiX1AQHPr9YB5gLhk8AvqCtUFp9V3esTBZDbWxFP
W9DGNGZKY051qu7bUnyhYNrS6eomMNX1AgG+W51B7YhDSBvI6F5osYMwUWO5wQQpgsCudrXiDUik
5TYQOZSx8ZInia0/TDELOE9GSJscJ2e7MQ3NU+20aDE006aoRt3nmWcW7ttXkcWHDlHNslbfW1PA
I9Zuto8bjxXNzpf1agN2hsY4nratE4qUW8/KdEtaFCK9v4r+mm8FQc+OSln8uBwsN6p7Dph5y67W
CtNBqGXyDR93Tu0UBzoAzwjcQtZohhbcGum4DuCLj/j5wghzQKKIA9xVlxOySYytjDlXU90we1VG
4KoZSXBwQ1rB1KzKQjckiujFut0dm8lrncNlDJ4fjQvlQ+q536ncgv+oW7O9c8W1nOrZqnpJEriv
OMPMKamtqHP55+vx3cZrmWlYnzN0sfZXsprm0OpVonP+Sx6Xg489IRV9x6NMhGjaDLGrxqwa+F1q
GxqY3Xr+gIdLK8UE+/9uorgA4NCEdpqrN4nsrhHs9d+pxhVAd9Gn4+AnMnhZi+8M6nw3nHXegKgd
WxwwGyeDnKEHoYAzchuRkH2EeKPIGuqwfEDwzjSCD49die2gniydfBL4dGfk9wI7ZrdDKEvAPtZs
glIXQ/6NwXba3M2coZNJYpFiH1Q+BErVznOBiSILuEvBIlFTKJzMXusUAnq9MFoFhU6gBJFGhX8d
r0huPScNEGVWHOljHdj2Ymvv6nd0Fhrki7W03rJ4WFbsNhKxijGHrpS9QLQgYk49CwKkscjszLf1
2FzG7zJcIGNqjaDWEIRe14H/ZPLfpKbbRiu9VY4k5p0ZCbBYSQUkcfGAIfVj6E/AzZ7HCbUfwFeD
/8cmDQLebfbuwreohvT9LK/O5eEWPXAOYrd7i9oj1fYPjdLniljP4VornqJLo4wLq0ZiY3W5o3A8
i8hz3h1KShuANFkXfS5Ik6TTvtC+teUzMgoMao0FjQcQ6aWHnvQEn+NzY16YibRPAWUBcWPsO00d
ntw1OrngefQyPQtH3aWzhj42RwX4NFX7e1ZE6J9eg1F2C1lFgHYQgEykexNHm8EUWL01/iDWP9hm
U0mRX87e92Zam0Eej2aB43SD2xmjaRMzLuAdKO637bSV3B4U/+eR0lXL/gMb5laZUqtRn9k544Xn
+uuWGW+4a9uVHuHZ5E6CpncSV74d51hBp4ObCu/kaPyuWb5ZFoC6EBDDJgje8gu7UP4FFCT/YZBo
UzHEH9CQwhl82szZBU3/UOiaBZKw9CJjZblDxS3MqC+hgi3nzcHGOAEteSLqU6AZnQhqN1UPPxfW
EgP4332OkX8yLSQqt7subLf7N1vUbujt4+l1Xnpb4juG1k9+2aHdqM2R6bU3Zuir56U1XR+aQ6AF
LvtDqVycjGSAe7MIIfvO1XejPu8+FDvBSewMm4AE5repY92ZHwDv6ZL12i8mOBxheoWHbbrYKeY6
t+wEIDu/NeUGL3EzBVjU4mGGUC8RJHec8qrsSa3ws44BjzwlBPB0YMraSjitYcnp20AxH35G1UM7
TTkKNuKlariOHAu0vVNot6waefDrh0tj2ie3ZSc5bdk6LtvMtUxle3mMB0jSuLo6axYvJYOosrlq
zjDGXLrpqzbCnB3QlvVPpv9sQvBO00s8WCyrLO7OZEsTJlFQIRAK8R0IV4UD8VJNyV5UgOdDmZT8
lgpl0uyTtLaFgo+ktSEMszcNMSKqDl//MQqVANx1boqEwvh/t7U5gWUUonkm9bHp8eFCMGEzVSGw
uaL1gl8TNMlWbTTK75hZ6CA4PWGr5RDY63i5NfxjLf+pr6BBuCIDjq4JaE92zm++rhpkXE34mOAG
1RVNzKxRJmnuwsDr7lTw82WhLp1T8Mf03lyPodFEkAjQoyPGcNWzMmSV7uO0SXcXLaPPobvwEA/i
EZ1OGXgD+pnXNkLTT991MUfaY6r27IJYsT6e8SIRhzP8ZMLp8IAMsQnY2309vkF2PIq1L1IGHkXR
mcbVvhKz+ShqxFGrwpX5UBtDqaQF/eQx1I088j93REyEQBG7eFGqHDKKLi67TWN6yz5Gx3hmj2IK
iSP5mwaxb/2XJ9UAGgsanzSSsWUWRIDNh+YgdFmrRxH2ZsOH4temdH05vCX0CXwZgyva3IfTVMvT
PPNOqvHEG2g/cJcZA7q+kFQbOP2vbkfImWYmwt7yHZECYqzqs0zjzYrukJDqG6AoIRJQ8s0Oy/ok
6oXqFguurq4hnIlm9JedjtUGsFoVxwJvi/hNtuTtKLDUPourgMixXo55PsCTGp4i5R404rfUZEj2
LSOxHrFOHKm7Lsx1uaZdIZLyKB9jDjvRpE7NBClEX/XUIWOMlGOIXMGbLz7+gZcwOLgpU/iG1XHT
SIbkni/6IEUyJwBdF9sDILetm63PRQ8zc802MH/lz0pueeDRF57POE1WU0cvvlo4J8bewFf5WwiQ
Va3PPEeF/3qn4buXG3CnRx4n4s3ccgaPQppf2x1HcxTqdEO8mE81OTb+Q1Heu46T8ckb2CKTHYEP
zRmxJ5oCMmXvaJSEiPhveo81bbdJe1vuE53/hP+enj+bnwJa73mjkPzwi/LILVqIFN8pl/IP7IXp
3exSYBEht502GTqCx8H+WXb+LsqPK8fk5XarjohUorc8zAZfQloUaCzqAePpR2OQ9kb8NLBK91je
2i8/AH6rv+W5Q9i1Hv4AJIJ8z/5396TpZWPAdMDvdtkoBle+kdJyjvrgeTkpo59eBvdqGP2B4XY+
K20zlcW8s3YqUgmmHd/rWt1I57PaxEc9NqIVjYMMvN24x/Qp9O7B+haAM6CO+PWWHgO+syvaRRJc
jMuL7qsFBXgGw18CFT2KUpIH+8o5eespMucO+y5p4pyYz/PWYJPz0hgbetRsANdtYgyJJaFT8aZ5
QWifMaRBJnjCHHZHpk1JvwRo25BxDb9evONH/qVHUHmhCh0e3rsezlCw2avCvglEMveVSEFSh2Sf
23Rfsl9wCQaYWCmUBDi6LhRPQB0hi8E+urcrawMgC5OnHOtgGz63BMIlND+VjncSEll0fyG6SyFP
JRj0jh/sys3X4rd1fYXn6COvzjVC8Xv/i9YIGN45G5HkGHUCbOD9sBmSb5p1anuXr5OstDd0A8Fz
6x2zmPDZfHS/eD9snoXkitZOt1P5HDPjMeAFvkjr3mFLBF/uqWV0sYviBh3aTTI0iLpubG0FOX8l
Nb8KtGYnRqV4WGcDVbKJM0yZxcx74r/yj1AjrNNiG1Br1ljF/4db5FUknDm5jdAIuwKvRDKYtjrM
EuBjiBm0qlUdauwzJSzzGpPXbVaSKhMYzkq9pahVfDVBq7LIgwymlHVhvEJ8o6uFhq4jOLBIgJ/L
a6jXidU6jdAwR0C5vaop3K1CRL4SSg8xSBQm9rSrdgujz2RIMv4r+Ah1kSX3dXia+WsF1jhscz8U
9tHDZoNcvuJ83/lBmD3zQAs2bPUy9m0ZRWee8A6rMe4DwY0CebwhFsDNLIAs7bCaku9vG5l/D64Z
7pEASRccmXyLzCrMjiZpY3v6rv3MeJmTnLtCFTqSp1vToPyjOLtq4KXJpEeaasPrjl9JRJtmN59s
xp1cGWzQMZsL+1Mf31GdVdmG5pr+30G3sjSMqwVhyk37Tu2XGx9Mb6tfk2f9Y1Y1h6+VLeULamTs
bDCe9xXnl0uQzzIh9FoVMcspuXCLtTJIECk+FXogrBJGjakkDrNk6JsT+FOoVe6umCnQ8HCeRt7Z
P187IAUAkpkYjYEukGCWdZe2gdWrSTMogmWzbSncA44qrSuHVj4aB8whjiy6zV/VpnexvU4o6in/
lnmsj09hboB5UJJZ5Z8M6DxwK4pr/ugrkFUMRE/OKw1dD0LDOwvDvnaSwRnci+UFmw3pSMZQmkIk
enQ4FG0KcYHzjPniEsJ06JeTFx7vteOok0aXMyF2S1RQj3UgNBt1Lx2YyTqJGAViNm3cadJcdT3B
tvZZjVadp4TX/pVGwKqun/Qp8y4eGkmwqO4UfIQ2iTPdPYEOwzuRJLT0LDJHi6doIkQfVLRume0W
SXm0SVgct5O4fwqgRDux9fpxaE3VIsgmOqqsm8HOLzQRJyOR+UyLeGP/+WXFOdkCa/1j4wrfk0aO
+WRc8kmd8MWqYO+UrJr12KmTu1XIWa1JQFXT+x4cJm9cltus8Ji2ZjvzgKp9GV0O9XkXtRndpqqA
NQHk1wJP/zkfV5YpQXab6JTYrOAQvsltmOOvgzwsn75ma7G7DdSKOjFwfqKwz4Da3AOpxQA6aBkP
5emAowMAMh68BJdzUADoIDP8TrHjnALRmV1hs/k53m3VVzg9BRoU3AvL01+E7hJbPthtX/zwTV/d
I5t89mvvMhUHxMuUJJsiJbbV/R5R1w9kP4RnI3gyCpVL+Y2By2EZAjPp7qpynR2oaeb3zJtcGFS+
zQDfK43XMdaob+1+yAiyOnc4kaM3FJ4yXfXjKiYTUc28IoEHxXoUO7nK4oSqqHPRcPoLbATdNcId
n2fFFyGzLJU7lzYEohqegXvOJX4outtRAMo9iRfmgDrzebnZj98Rrr4jZOPXQNrQQNCwN5ONU7dd
n9MzAPC81fr7lewVYc3+dsMm3V6AcdxIvaGrJO9i3h8pU1C8Ly+EiWy37wUADW8UBgyoSjo/0tye
xTYDYhhmcx8hcVFIVg5SnYgWqqyC5eTXBfI75ah8eu5hAtFxyHyhX4PF17/LVwiUCY02BB+N0eJL
GY/7HVs2f12ckDzkASp1Gy0FXrsStiFNNU683kzBhkHAdOQhDV1o/d727888+0qejNajm3ad+Aqz
RPl7z4oNrEC74a4Lgnk6GI58mKKh9g9JbZx2Z8y4ZxFfIfRhgxS8S6BY55v27bvQ/44bVsYL7J8Q
LhxgqCT0TdMmQZsiTcT2g1bSluS2bK32fUGFOlSzU1sX+UsRHZOf0h48IwrxT74wBVrPxCxjzOyQ
VQQ1TsX2gEPkIPHVg6BmFDJ2OxdU1/S4Z4OIomvtrDu5tyu/2TrRHvQuLicKaT9gh9sNRHs363dS
nzhxtHRlQR0/QY09YqwuCVX1yuAGiBajBl4EZm9898Ctc6RdemfxkPJlIjnSwR1ZekhVGASpCm9D
70WjT3CRqRHG/lOG0IPL0kP2Yu8m3JLlu/19SZFQKZIXwEeuOeNle2KoysCbSjk5L0Ht2YGDusID
bFRyPGulrDXcA1VCWkyxTApp10o856genJsMPVlhxKdM4HruHnRDEFONwRzJDRk62h0PuDPfKUui
GWWb3UhhlxQ/5cSQY9xZdOkMIwgSa8AB/AuiIzquSXsj8Gq5gdgY7k7uhiqjUKnB3FnxM8TdbESK
8iCGb6vH6VAnxJx2g8HuKlC/OaC96vxETSFWKfc+eK/0DIPW3KlWJklnwzWo+F/egTBBeOob6Gep
evCSOhG+8zgYqGWJzUIMgtNyrmwcZyXX/FETOPG6PxSSYNNwM4ZSpcvbmw+qgX7d/Ye+NmB0fzy0
U0xg5n9x4qWabVPqrlpjKmwyVuG7h2duWGVy1bTkzTeb2EjK9WhnbFuUx9jGzOrHqqtYPUvpG1gA
/wWw8Zz61SWlih6/tok0TFjKFZz5hrQ9DAETwtnJGlJgQn8IVxLy0FEGijONBwmUSWjMnKJISHnv
nMJIUw8WFXdc7iN+KRslCfCvHomIqjb+3+ki4r7gmTQEsZNLUwd600J1+gFCG3H8IvwI9OWmq+S7
dbWiVpjoyNdR7TI7GrRlgF9VwxdjoIwsEjVxSnIvdbxQpKl6tnm2VJ4WzEyS3ojStk/Ci1K97WCb
gNCzOH06H3Ao7BwWor+7cNT1kX4LT/MlNGiAHWyKDDMuOqVkfPszQOvyeEAVN7um7usSNr5VgcOz
xvm6JbSdBRrXE5D2GStF5Qa12fIlGsIp9Wr+okyJMUIXzoxBtuZf4/qQZalKgh0GXF5/LTFkokkV
4VGrFUcnoJfhEzVHKkcQnk6q2noBJ1FtmTuw/hVN/q9zC835FBzNG+qWY484O2eESbl2fUCT5ANa
gOKxqPByYWmLz8aycey7mnJZNipQyDDB5bP+Nj6zrdu1XElxlzaRJ8PuywhjTinPHp6O9AO186o+
J3oNEv9c8w1+DGe3Avi38xWQ9BFIxPbbK0FcUra0z87NUK6lgIfRqj1FrKEiGzpF5BK0s4Xfa67u
jr0apHUcCXgbgglY5hptCTEFqenlnCtcXEXqEvL6nlW6PBV0xUcXc5u8xpDduzTcAhaHhZj50i87
I/O8Td5GgW3P/yZntHQ/ALA9jjSc2Q+0TJTTgUMr4Occ2TlINWmBkkmcMx8NsDXBibXmNyzkad3Q
WISWBzviqvSQkjVSAr6tC95gQDULM8lueiQYML77aaRb0zSNEjkDyYkZQPUN/gEXofKHtQqxttIV
D4k1jJMDDFs25rBbG/134ERKxa6ON3z6KwFutTnQLDNeNb3BkcEkLwoQMb9FWNvG4iXKMMNWPrWb
PAsraIYxiKMRP0TJ2o+YGdggT3xBlmQfKYaanH6kRXLSAUfOF5PVnOwIMzNY3foVu+qEOkc3ztlQ
n9cTBLRxQg+65F0h/bD29cI9FkSzvAgbIxAm2IWjD728dGFxiDiBEwEbkiXiCrwiOoKz7mFFHAqP
ohLyGTQxCJtgp9Lj4rgSz2UgrVOrpze9uNUiM3GEio2vCH8JW/r2iCJGw17igZNzi4v/OM/kFkBO
vW0ffVUfTcrbMlLZUwp4/r9NHSqe7SrDPdgz+IYSlRqiCH2ZhuApTj0PWsRwCMbdLmSVnzvz+E6E
wetrff68rKeS3b6nuSZUYxktmyk4q3WYuskLo/d84DmK77MF8ZmJFbqA2acp5g6zSjPYXMUaalo2
T2f7OtemalfmITLeAFE1/OP8zoxw8k+2Kdv+8kpmpJRf2O/uIAi9NCD2XlmcOGeS57/O3rwROvNS
TEVOpK7kmwtR//PfN7XQvoyAsTgcHt4zc2ZcUaHcWKb8PDJkUzaHI0Fo8XJ0XDEi3jD8+lU7Laak
rZ+lskelSLD0ZTFs+IHQDjhP+A/LfFK4eyNMLrXgnOianmq1UrgcWmHaE/6cjzJUwHiwDs6StKsI
rEz5piucn4EpSIr2DvedcuUPAq9/+B6gRj7LoIdpYgzN11+MVTuMsDs4iIzyuraECTIzAUgzFHkk
pihUZ8cDlb50kQ2HBLY5X2t1FId4uz/Tn5x02mYjFJUUQFbeNUT8kLjlEnUkuOWjCocG4xd3qXsG
kV0fbLdod/f76DRQverPy9k1flIzz0NP980TGijrjn3YQKXvS4BG1w2871Ohc9ss3j+S2pxCMGwP
lKVxbygZ4cN1Xc82Z/1cMg5XFlistYkpIijzlkXx4KAxgyZ5c3oLBm6IF5iJkh/1Xfq/FV7uLTMZ
F3vb8NWLekgQ3rUojN1zaqa3ljzlW7VBFbERUOEjXviR+GakCB72JTUn945MC30auu5X+rGUxtm2
7VLL4tQJ2i/C2E2TaATfjtqrB3Xde4qKZNgBt9IPBNY5qwYnVV1MC/uovjc6LrL+1XGo9ZXZ3p65
WPUU+TERKGVl3Waih7eiT8/0VaQclUz6oR9H6mAosTomi50pCYoxFYoYRRT7bp3E0s+iE1iYAxVl
tViwPMlU9XMCx4aZPscol9MsCa3uqnW4rS0DOKkYIBlzNpUzL/GHl0Z5S2ZYOjNsMe3VDQAlvTB1
WWhKgKLbh9A7xlmxR5Kun1x/ryVcrCS7ITVY6+o+ct6USpxQY+FHp9J2qQnOn1dSe+jKj+2n/yQe
/Z2qQtO+MImeLUYk5u1t5pfjIfQjITtnNjDOMSzYGWO9B38aFMqb0PgEX4JjT4qUPxQR50UR6fhh
4DQcnpJr31NO0gNqDX6ixedEPreOVE4BumHGXyHf6S59vKc2JJbXc6QPto3+l3WxmQTs8ELTf4gl
w9002wp2JTsRlfTZiik4ZSDGzo9zeVfiGGyojfMB3BZjSyP6aIT1KP8BLB9hn5bLIthH0GWeJN8E
MzH1RLzxsQPuiyYXnJu9qkCJtY6Q5E1fGfFsL24ZCJSP0flvDIIFzPnm5cxWZ0nY7cfeczJNCq5S
5UUH9bhQ5cQro1SlBgUjKcZhwnwzklAhw6/Ux4572Uzd+2mf73GTfcRO3LBUnzycn9SN07b2jsMa
6fZqh5pzvnrjIJHaenQsFl05vUbdu/yrwmOnKeF9ceN47bNEPCMN5jQaRM48tqBbOE59ccjUQSp8
XfJyoNvRAdvtBZflVv3edS0JqHNA8oOnNFUzp8Te9Ls3Mz2aSojbJ38zSH3iR6xVzDtasU0KIpEZ
d0I0XwEIUq/MEX+PBmfGfz6f1uwC/hdK3Ke8YoWRJrNK3YWISQpuzBwnczd6Ar8fuxylm/WvyLFh
puIuoqc0oloUSUVc2HYSbJ5DWA0PwdwjbMIoT3y/Jp1HZXbtXe0ysXqXcvUnBXZiLBojx7MrzsMG
/H8rtzG2Grckm757GSCouVIEJhKCBrzLyljG+24lJnBmbKLqTy4rdnGvwNTY75Q/FPaFMlx48ff8
FzjhRcyMOJIb9xGLlSQXp8+L+x5q283E+Mjne9Oho/icZtV722qIA79ax1pMWVgaL26pXrE24zj6
2/ozFgc0qpXy7z4AkLf3kGSa1mJTQzNz/KzsaCgDHE8jq9aR1zTrKBG3cmdrNMAQTB7suUKn6jGM
ur0Q5A3U2GBznEPQ7Nw/mfXGHquJeGbjZjoiREKXshZ+EhcJjuDCaFSaST6rVgdeUDSgbb99P50K
VnlQsoUY1rLbOSdcDQAf1a1NoLKBzf5U8sGGFGkPvfTMzP4TFAuDQEIgP5+WRY2Bo4ya2tK+l108
uKSbs3etuWDeOch4uNfN5DEJt3VvW/ug4aOFRE9fR4H11Auf8+MBjpdIxV75qJOAIiwJ99th7OJw
YrHBB1V+kNyMvuEL6gCvMSQO3pnd/IABG9EnDre1BVfIDOQhVmjq04fJtIdYdoxgrLadHpJbIh+d
nyG+JeEXSHZuxWiYt5anw1JlSV1IUMYbj7yxbG2c2KwTM1+dnfS2R6YP/4VdgkeDpxENdTYb2LOt
cQ0y1PsWmuzuhMIbRD2MO74MNoaZkvW/tGM1tntuqcArHI52Ivxo7YQAvAZcaebm0tECJMvx0MnU
oLpi3RK0MSa5wSucjFt8OACCEgYhqvRH8V5+Bn90eZuo3k+oZrXIF69Wra8mzfuDiLAANi11yDI2
FfljUuRV1hEdfFuhQ1dGIwpmTcQxby1+AMWwNUTgUDKMCJ086LC0T0kDR6ftLumRxecsUlUyC7Nl
0S0W5OtxGX6y2GktmaPFdRUjs8t8h0DsdZ+qhZLyvnM+ReEj71zu9rN9I+Gkc++6kU7TWmUOElsT
lho4zI2nk0jh6oCS6LO7iDFzcTFS6FZzrAlhP4TRa8an+1RhbROX0j6OOCtDbDuurmkixXpn7Ya3
p73HdQYuu9xm/gphE0WAl/y224maxgNkQLNUIyBMcAHs5EtoVAZ0BklHvXEBqAIJo2Wxcf2p50iN
iknhcJsHnDE40wS8uK/23/XU7ixKmBN5W8HO/4lVFTGjZnf1sbVn04xWG5ef5aG8i03KH/1Ft+0P
WMQ+4f4HC28qDPhSiNWE2DSZxQ1AN9fWGQooJ0gVBUdFzAr2chWefw6+dgAtjOjis+HALoKUB72F
scwiP8AL4mSd2Z7hI96AXQOx4nDMrm3hJH8CLO+XzMc/zdte0Q7C0BjTUT67s3j2vYMYc6zn03uR
CvuG1hJ0vDZgx8knfHQHs90Qo+tI9/i7BUhXEAtneni3lX7tB10yp4LIxEDO9l0grSq2E+VTj4+J
ZCOUk5suRQb8WthRXXf6HnMhUIrdNMm3eBag5ZECM18wMX7GT/rw7B28n8ks9PjdQbLAMH65Zd3R
1UyFQ2z6igltmVkzv4hKfvBL1MDPv1+SPQSa0QcNeZzAfA/3VQi3DhsfPJrcuoCeYdmctccIC2AQ
0o+3u27EHDDZrTYrC/OxRssEx9NT5Rm5HiOpGT+odBDZcV+QFAvUzdOyp/etSGvQwbJyk7Z+JpnB
+t5RukosbsL9XRi4BR1jZ6Z7P47LakaMYS9LGiMVDjSRFszf4T68nOfvRSYIk71wAYWT+HulC8Rq
vaVB7oNfh6aUNcOy7mYZFzVEhlaJMUItDW9PbO8CY4M/XJoCHb3zp+yc/MoxeQGws/38e1PI2bxl
ReMwRjKnQiAvZSn8lm3JTaqFOLd+baJmGSxjUFnJt011hrK7Oahw6o4nwqlUBwllX3E1OBJlUxoD
0xlYtpYG0YSBcgjPklz/an+X72Mk1NGLVoPmPo1DD+Iqf3biR/Dei8m97HIHhF9UDVBVKDu+EBHS
wU5e6beScRjQwNOKnLDCAG440eAsdQhndORu0G+bpCkwlwXjxJ7+nLyJ/2V4lLmbU+QQTG1AC/kX
3F2U/MXB+kN6cnKBGGtrIBZqLO7pBCa7mEcKjvdiF1zPKJ/tIA3qGA2xUkV7sglM3fZBq60X1r2B
0cQ7JpItsbbeJbbFu59A1sOuwAOhx1QKR42CwmO1bMFR/8+xulb6VQJrLi8cQYRJUhdWPTLqlh6b
pDBqP9F1E8EGdm+nOUUq4X8lNExtlgK85sSyVpOXWGClxpS2+xYt79hkirMsb1spwVdyXD6KHgE2
Wg6nSnPPUx3u02R+KcL8nErwPutqML3OQRMWeEgFJEy4g5U023LXGysl9B5YxwStV9Tzrv+sY/al
mojEazmxrJwt5jkySCcx+XaROTfRyD+uDkYcwkb+cFRd+G/TmMSyAQAYebtFuqdZ0yqlmpxJIlrF
XcCfQNKhbkxNefPmoNpqQBaF9TFPy7BN53EO5aij3BRhRHlu+0O4ng6ue86E6q8ayX6tuRP1oAF7
6ulbMOKcjWv3+4IGekRBARwqC1bF5xSNi7i98V74hzojLR3CMzXZWWZUul+HnWBlN0zvR6EIQDwG
yR1lLbglqlbdWK19xuDHC7y7WxqIRj6uDRojE1/UBrBRLNx/S1BoJDvBHCCykH7hXOgXBPk9WatD
s5Q95nMbyVQydcSjHotylsN47wVWBRK8YIMQaIYbPWGQ0xwyP5FZz4wi1R/9eE5fccFVNMx3Fp3W
qEeAl8+1fl28eVdfo3uedUO2r4VE3TIRqSCEIm5Zvm6Jb4f5S05JqHAus/8Yh+dqN9fvRNTnolsr
G6lRCzBhz719H2nZfv1Z5AaZZpVl4YL5vPB6ZKB0kGNg9S/FEG4CYUR4q+GPiZwdPjsW5m9L7Dtl
dGn+s+CpBZBWTLgS44xSdoJhbD2alxp9+yZ/DlnxWHTw55Qov5Zg925WKlAFxeL8zYG2lnJ802+x
Ba77WP1nSFfPPqCpjSlELqOVKLuliGyMVCWL4tQWp1I0+Dca1CYTXi2no0kDhSmIv6cnxJdGYnwf
WXKX1ui5VYT7uVC4B2jRfQphcpkDU1mEtv/82I2YE8xf4yCX2cJurwx1TcJP54TouYMcjiewKAZ0
Mpv6ObkCqW8jLZwkYo7p41H5aWgTwSzCrJlkCtiMCDX64bOH19UyOSkN7QmsBjk2Oug2frq7t/o1
h4/YhqLolpnk4BM0aOlmBrS/b+iF8FoaZZilu1qwNHCIYgNW1xJYHlnibDbvqc5QHQcAZ1fHP3yv
V5FSgUfPTi2G53/aB4Bf23GgjUUWMqh+k/9SdhgbJ4Hm45dfjINnRiwLrGI2xq2Pp8eCUCZP++T0
oPsqAeqZ389OtkhHnkBYXYDW//sRalwnA28Ry2duGgaQK1HeaaTImtyFvUsRo8mxz/u8Q/VWu30c
Pw1vhLgVhkAZbQerazQY8rwr8DHxJn3xpUtyjr97M7p4xnvUsUL2hojUDYjmYefbuIR1/RLvx4CV
ide0FQ7NBQ4EaDw57Mvy4OuhkzBkC24eQPyduDqZ2ITh7yiqT0zzdsKSomEK+sBCYSdyoxrvP0QQ
1EYKBSQqIyvl/6SBbO1b/PC29JFblYURGTv7RF8J1i7eqf0Q1GmglmbzRRIOsxkEEZQ5ePKFkQlh
02cpiwzPQWLI2gLfISzum1SX6YLaMX/s8FIQDlEwPwPHmOusJhEHlNyyvndri+bobL+s3hiUC+kC
deV95/AFcAk0rSwXDRlPEMFkV786NlSNNqJ2tNRC7y0Mqt9gGJCzll+XZI0KF6k4XvAeVYmZkuJr
/KexslXxO4XHz3z+T4Pil9XLl7rd+Me6SU2uFP/z5Dagt4x/XtJ3h+1Sza+YNf49ijsKZvyIW6l0
jdy1otKyz4V4USQtQBtHG2fxjrWGKmzpuHBBdNRaGQz6qL1OJtRGEfn2ltE1VKrQvSWhU3UDcKA/
i4ED21mMXf7DWZ7aFikEdkrggEICs6iV5jL5KWOaSgSauDCmWMLoAzpbr1y5Q8UKL6FCq1Uc72Xg
SF5vQSaLzmLouvaNdAV8cDVFX3pwYuh0eVVfsRDPGPnfCkeaebkH0wSwgTh7+uZB8zfD+L1SXs/I
1XfeGT8/iSrYu5pDCsKcs9gvdc7dhlLPqIqf57796QrK8EZuCaaatja/7FqudoUdJ0dRUQjtfEVr
SgxLxPL1UVd4VBQprF11vJJSNCuJlbVMqEppW0LOC4wJu1lZVZ9CivHJcK66uP1+i7EZAOmKiR5h
3eoFsGEZLsFgoOSi2ErcNBecugbp3IB8LmO5+/kgawB/gEGOEC1YQxc5vWhEEgKm70Os42Q0z7/E
umqGW7hovjfNaceL0h7+DAw5Lk9aPZtSBCx7SYyn7uLZ/MVWbvNPT07YCuCO8tUp9pBbHjBJKJ4O
M14th5Xi3XxFHwqgBHAtPs05au2L9Kc5camBavBqOcxoQ2GjwFF+vV9Rnovq5HmALpfm3sh2WsgS
igPciEgznQLVi4+b3AeUP3+YZ7pihVZxXBvne95/YBAir8SY6vH5SCkHwztHYOcL5kTWVffnR7Y4
UJ7GGcrlJ8+o4cj4S8BQ0UOKgNr1E9t9Lu6rg9CqEVzneamFSKF4Xv8Y1KurW+Ii6S6alVf9ZqiB
idPGTyFRvdtOFKUakJ5RL92s1aUXVkNsw9jLvufklVYAOkbP3Luu+tvR90XN8uaEb00fCi+wFkU9
+JRZvtni+SqH/Z6/hC8xPOoyrw5O3kqqfzb9T8MKDIVozqMM48SgSxDmdE6506JKLdABcOc8L6Nm
G9nGv9g5BROTyVxW7fk7yrv6P1ShLVWi+2Bj26QYF6MmuMqKXuoLKd1uZ5ziXrb7z5oyJ7ltUHLY
4ME42PJr2qTo/sT95n2R52IbnkImDvaVxjemHeY9CTZuiZjInk8rXldgljClkYWz+8prtsMALoew
EHXGXXLyocH6VdEH2iyxjdHWGnNATL/us6McUFClJvudtsw3cfHMqnMhjjyg4WAiLBGM8DVupBh+
lDoL2ZhjZLA65h0JRkA1xjhOHnXbCx7h5zDUUPakei0SREcynlR3XBmx+ObSq9E2Uyp1pTo773jp
Fz+VI8k517ag5eLtwjZSeYcETKU8k3cZY0/+f2cSN8pvpGziXCKAzjvvD+5GwfZf/zRDXyOoTBc/
Hv9MIlDTLhCe3bphSor4rMhhURLpjOiSgOSXcjRalL7ODdUrGVAX3Vm1QbfyIFiCN1soM+DC0qGE
aoFRQPSN2dYpJ+XKdT1tqS2JiKaPYKZf7H3GaE94CLCdt0qLc/l1jwTWhZAoLQuE9dhj/nGzX2Un
ameRbmwemyv3DKWCKghwohb3A88+gsMyGXAOalRz67HmJIaxmKhe64aYlK0QkuEZ5IF1p4qNEpKI
8I5ZvPmSg26c+jDvAE5V+GzE+HA7xv5DCPxdABwbD6HP1TLJ+dMLHbDiJvGRKSqK7Sm9Yi8/Oa3/
ECwKRZrEvNyK1nXnCoHq2zDnHUHN3MyOz36038ZKF1tjB6cSaE2SKfHQHHAgr7NYPrRj5GPLKHss
CPA0de8cLBQ9byC+FkxgwllbL9VVpkvcYSZwkJD1GLIjoCimsva9evPFBlZT8Z2eF7u2vRCo5mfi
2njodN2gDPgdwg8dxSdwxdeFOdzvHnMOOQTH4J6OtfoRF6gSvZ8AoZYrOUhSf4hx2LqjX3DuMh+r
zmKrLeY0RbDhnZl3qYrEibInsM/OMX324wvLFPcHqyv0hEf21YvjWiyeq5PDCEgSvYE5jB0dfByo
u4ykB6a3HPeXUr0n8Wz3xLVxoKg72wSmk6ULm32y2bW8LjbQFJ/aV/zRt+8lOpyhXsHkH0Hv8/4/
/JdFUEHE7WWhpFFaO1xO8L6oBFuElnH/93cg79UWJ9MdWaABNKudtjp5ayhnHWKbOpFdjdoBOjrX
AIKaoNqDHJ6S9k1MHaE6uCCW7/fRZeGhVOFeMgL9PCWyLE0tfEK2FZW0pXrOESDd8Cl7J/4Ekyns
x111Tl+lXafszVeXQ2USeiXLnhNT8LFckHeRHTkmoIp4NuLuWJOdOyTytd2XK8Yor4hh/dyg+9Yx
mj3dJvRwiD3L7MD8zFADT9oL09hM+wilXlK1V4j+A5xzJQn55vgNRaANHuP+uIK9JUlAd/uk5p0B
dhUppzGvxWtUV7SC15I+f8b3QCHh16PFSZuz/Vfo7ebkaosgoeqnuoZNMAgluQ4EIlqTCeXxfxoj
P3G56tbCnxYLt11oBtcvLR6++7R/g1fP5JctjZlPwRyjS5PLu5FgIlMPXljWvt3kzt1ULw4XfbC/
bh1bbemHlDCVUIOcg6em/m85L4EoxJWP7EI0ZmEt8JYs647z5hsrZJYPTpxCldlnyCYt6ZE5Sffp
X5Ss1CAfovEisSFMZt1r6iTa/272VY6+P5Fah2R4QeFhPln8PeFTbSTAljJL2+vMQnRHLPjHttZ6
t/ZENhkaSy7ipbBOgsW+SsbJBenlj3IH5UR5DOxI++kRbvpVzDuFcJxqzlj5YKi7dpqRGDGtRadY
ndF2b/vX9b5IC8i3B1R9pOz8aFM0nzGXHWPL+Cj/lDLL4iUEhwTmKkeU4+p+e6qbFOy1JYd/1+W0
n1FXN5iFFqR6G6BOK8BzjZuJyIn/O2i/L5eeU76jW0qmYEpJKK4DGoKYqdC9Yv8EnQoZp0gIseAi
qSXdmCKLkOLspHuz6EQaDGtijE5zeC/4Vs12NbYz82UZseOxyq8naXBy9FqWqzhFK9RYaUgYR6yq
M/79K45l78x1ch2hxxYuQLeoWqrRwII+2UHASiJfYmcDtA1PFJbejEeZVEilQl8Xh/P+W/vtlQHR
vwvsdC+BWeUvkEdj6mFANbroh0iQazfaPHfkZTD+bWZn+sZey8rAtUGGj3fjhkspDVR/CeERt+qJ
+TEZbDQG+wNJqE8Td4k4Ju8s4TLIGUVxztdrNUOpF6ydSYmGy0oRvtLkIw1oJbMayX5PzFFdQioG
ieS4cb6xkprmsWIV/DEjjGLPc+b5E4YF9Ul8mJC605pVKM7S74KPeb0wLOqc/j1binLgEozUjIeQ
LjZ7syQJS26Kn4Mf/KuocKTE1HnpS1l2s1wsUYYmF2S0GCehFwvPA3/DwFLa5lAcXuD06K6AhozR
YqPTsQ2UKqqHmAhbhPvvw71h9xf6sawR6WAVv5ivqCcYjFvN/ol6ueD3iAM1hv09A8ekWqvpa6z4
otemMOnliMyy6Y6YjkAq+8lKpjQVUfLplm9ziTJSJfS19SpAOKpxs1vL0u6s72Xnzr2M385l6gyW
3Lz33oB77wmiy7SCK/5sUVZ8W+slK/LuyGmFw4XFIRg0mKEC6Bj+64Z1RzT89gujDSBa26rYgZAP
vPOEvm323IHclPVM3EZZrNrVi09zaIj4wooAnv0TmEyP76yrPjit/S+z8SQZQFtm+lc08vI/1+KI
LP1g2SM1Gmli0ZPXrNhQ62FOur+6WaemwHTL8qo+BQW9Eex9uxF8+GtBQhH/1MRH4JcUEKFW7NxU
LLup/1BLSG3YdcnYlaGStWXw63AEyiwZezLutvA/zsQ1Ep07Fb5xuYWhsQaFmFMrFanA31Pvroej
I5sIG0zd0+VK18TczYrKrCkJl1ou2Ok5BqjVhpeOWqYNQiPNJzV0N7UZi8WL+uzElCHEC5+VicfH
pEkK7dKM5jWh5pL/o7CChQK+EtJbZufZNlySa3fKWo3ICtkVsKwWjdhCqL3leau/K7GIbd9ZuIov
qDQ5KF9zIdX65Vnr2+8RPLl4mr2HgzHMq23N1/DNUuGp2jMmnuUH/J8AWGcjHD0GbfIfQkO2n832
e/hDaaEGmUm9XErzmT4+eK9bxEwXomkph//hp8M9pq6ac4yOltFTPWX3fmt7lHHUu2snU1p2KdtW
YG6LmS7KzJ/Z5sPj3EpmKeyiSrAHx5gCw1r6fJZII/Jsq8OXvtjt3tlWT9KlmTX9nmENctxauvOR
5pHrF+NJNV/GLbPwhQYNZJJL60irw60Zlhe/C+CHkNgxuqyRAGGt26TsguGRExlZCqATcshapHpV
0yFWtC2P9qNWR/b8YlYb1NsX3JLeyduVNqCXDpvROO5NJkqg6hvrSxd3BqV07JBVMQTv9jtFg+Dq
LkHlEb/j79PO6Y5SL9pCzRLSjPx+SVZ7PtJTMRR+jB2b2uG3b1XO6+7APli6AhkdQqVJN4Qj/ahr
S3OOS9tY8X4MDLJpQiA+58fEtty5n2W4JxggwXq3CxDabeiWUyUzPSwtvyEKvgzwuNa3DwPCldnp
ZB9rK/LMtIJ24sTvU8MJUyfCC1wd78YRuzA1wazNa/NEme/HyGRMgZHOXoXmI6IathOlO9MMnjQQ
+ziPUTHl85fk7XOm161RbwaOtpSqDyFAYAwN6JHkB0gLYmAWTypHIjirGMK5DfRQ5D80b6mqdbwD
IxbC01Op+i41XZGUV4+4lUsZ29aO81Z5aT2kFVNSPTfhCaCKvdwD6/1fJ6+lhNnPV6bTCsEW+T2P
XQcKXTLomz75nLB4GliZt/CMum50R610LgOjVosHWvTSowtwdaZse2RiUI8k7icCYIKSlm2mlb2U
gUJlHzx1YjfHRUj2En//D6VlNlrtkUVWcbZUEcyk+3Z1A+UPfU3PSWcjJyrcLS7IygMeVR9kWKS4
honXprn/ZmVVP7L/lG/ojyvCyFBPh8dUaWdUCgofy5g3COP5IV42PbV5LA5ViS+SIUNyuVaqoMAZ
qxnH6SC0CvWqvnTw/mUDPrl8OIySEdJH8i16W+SQOAOoddtTzyYi5yqj0figftTEhOmViKERtsnT
4iYuXuMYMSvnIbnFbEW6C54Iz8tkzlJHSHLi8mo/ZLwx4YCUYClhpyQkfUDOoHy+x2GWh8xlFAJE
C7A+a+ccy3D+aUEh5dTljcefSwuIA+4Q5j2ZuYpgW6GvXe/HpRKaEIVzb8na925NJiTR0jLP88V0
3Y/gp+nQPV1us50N9CHkHVv9lfHN4LqEJkxvMK96endDXU22/X6vmCH4PJbZUoPMNz4KxMg7zDQn
D6CK2JrsZTrUmoBfILqH238qGlnXEwK9S2nrs6R6v7qNmVP/1aZm0Z37fXpn5WpUODWfThWvuTyz
BmneGbzaBskGdGDwywNaNeV8MrxOtWszv8qOG2DqBZkvTqZh0S3c00BwYiA1n3ynvvCch7s5sMcQ
Y0YX4+a4TdeKTxpeokKijusvyA4qgzCsoP9PR8G0ZnogOgVm6N5XAKp/KuVrMZ4qMqrwZyIae4Ps
lr4DgXAaKyIDtdSoWFVMECFvoga3/T+GFCYi3eRt0nuAJsw2JKdFaePDyOn2Dj8PTFJPv71W6FiG
wz8MQW1aWwYWmRPSChDVt6k/zg89REf0L1qDmguzv0ljrBVVlLK666HeHF4d07pLRJ6DmJDvts9R
ApMFNoeKWAqPqJeKdlmnQWqWlzbEJLByNxOR50+m6KQjMa4Favx0X2Z+mNkMuApyHGslfxrwByXP
Yi7nNnJ5IB0WA7UpXoUPAwSxKBNmRJeViTcBnGlv+/cqd2GiHNZ3LtFU/U76z13gamnIDn3kv63f
vr9fGUssAhUJDafDljaTKqQfqd2c08hVxump3S8P8gB+hTxXs4k0/VnrnSR5iVokwEG7JrJF7Hfs
Vs9c10+oosjyUHKD0wUIcvxUDH+0jNeQaHo6D3GjRVatHaGZ3eL3/G9WTjBWFB+QQ2cKWQRqLR6t
M8YF28dtArAXW/p9gzk+brDwdaiIaJLC+7cxMPhunPvlf3uzGsNqUZCSgrZpyOVSMO8DLcFMsorp
YcD1rHtjBNGwe3IGdn+kFyvrXgNSqdkaR7BnzaA4kPLwFHFmOhaU2BOX9BvjErSBKFKVthGQn6BP
UHCqaAhqi3ms57vqz0KJcuRwwH91nLamCHI5dW/0nwXWL5Ie1H5Yx0a2rHxqqPUuG3aDSN+MzH1H
ee2TeN23Bwj+Cw4YcTGEYnE1x8KjgQtjHaZB9Fn1v3aG8WGtOrHSW2rlQwG9BDtC52XfTtyDYfHp
Tcs6jRo0jMjoGvOQQ+qFMWso+WTxhvHhbKcMrOdaDqEjqZWNWL0ZhsQ9Bd1C84/jJA1rBH9EsUdp
K9R4qGWktPRkwVW8sYqXJcFNJqMU2ROamS03Jhorcu38mOyRH4qkpzZnQIMSQJzJYohLan+szYgE
DDoIwUStz6DY4pZFKygs8AKxKGp3MO29EBKqv+hX4ACFox0TCooxOd0r8MRfan0pMr/1MsmMDNho
K/JTYvZagzZuSBcNW7n+MbQ568H78rrx5QVABiAFyP0ShgFZoCCmEf882nX7lsiaLbbI4OfqxzEY
Dd5U1F6naS4ar3DoJw6w9vsQ4jjxlUSumC0W5YfYROgghT+SBow5KjDb/WZDl/sSFbHmFcrc8AQe
ia+hQ69lDL2RwobRQLS8JMm/vCl/p2fhEojD5bI549WBJCQqRyJlaL9RtANtOO5bRaSrh0kqwge6
P8Ulkyhwg1blHQ06wfkj5GxML4UKkDqHEz8c0T/IHqSP4/PqdKndPXBEw+WS1uqc83ciWFH7rGjT
MNGJNSCNMJIxCUyzT7kDk0y+GQivN75qcOPXtKtAIO+ifYFF6qd8QPXWYNlM25kKAo6gD/xWQu55
Du5SKTWN1cr01S0OnWJJ5MVtdepWssW8inhe+/y9MH20yJ56W6kcXV3WmB+Fesm1Zu8DW79Jy5j3
2Cd9F6nPJ65C/tLjXEW9fY+oOI9/1UdDDJKMSiNurhw0CMH9iKS8grezVn1d+GFgKlFJVLV16Iw7
XiO6Ft69G2XDwJszKBc8VwS6jcHIeMM/SLP+S1KdFekBvhnbPBAY4s+V6nVo73e4rotQGbJ5nycg
Y1I+rDHyJJvGgDPacLxg0cdBq9/mATMHzn/3isggoF63UupA8ON7YRQ+Bo7HmFf+LryAcuQzJuh8
M7oz6EPTE0VZNo+9TOI4wB67fv3KcG9SV8yMOsRhvU4KnCXG/DKccWno17gAmaTV2FyqDGtjx86Y
oGVmOFW03z35FERIc+aKwWiR5XKKlIgfFqsiVxb8Ti70EzWdzrjBMLoSWOF9CdkuZ1uCw24tLrDU
vPk9buad2S9UxUxAwvmnj6IefB7QOlhAL6q5kAICPCCP3fTvu+iQJ4EJRRjBRxdEdhlJvDUQIZSb
GAIQj9zST4KeCHQDa7NLMlR4IThirEyNNMYemRJwfwi/5TQU6M8htxkNpbzA1LZCmNaMxFm8DGlo
+9MDMXWsSUVhj48MbZnCMZstaUpopqD/KRjxjmoNEbAXvjPCoNlG8h8uZB11ufhHZ/5A8R4NzhsN
bWpQEa3mKvP/O9VJ4shHJxF0ggQzRkFEhpo4W5e9uzzMx0a9aKAabpRL/dWAJxgXuz7HTxt/5fLQ
FbaUx9T3e+7DGD+Exv9ecK4pxEHmmJ4uEyQcowzTrR5UVSl/8PUAhps/sP0yU92p6sllkhAsUebx
RLrMGBEgdNj3aoYnMjpZDFtdUlp+3diPK9fLI3enOzHACqpC85ZRVj7D4ofRaVKra8LET3pWQoVd
66P0ZBGYpZ4Ux5d0g9ehvF4CfEEH/x7epnlP/dCnyYuJKWSeshofFFEh5yztruOx/brbtT7wVkc5
CfiqMCvbHpniPzksOQN9AxICZeX2gehG3N3VyuOAdezxQpBLoqsyYcnruNJUGCVh9bDeRDxWMK0w
xK/DvxEjuy9sx4Ovkm2kgvm9uy94kFso6GgMPAIRVJtsCgt/lpupS/cVb+gPb95OCE29iNeKDYUv
xEKiIYItp0UMvtEh78as/v+ejR8y6IM0UW+mxoN1C1G68Jp/P3LSCac2oCS951rvUzYgCnrdhcKF
e2mV1sc8DkPJpqq/edrW/0I+bpg4V2oBZ6oiu179ASCP1u4GfziKZ/Rj9KKo8lZVaTLl5Vmveiq3
SUQAFYeGfMGTUvYozyJK45KbyPWUlkfZxg1NOmFkFN4dQj41Eigz5uaQNDdq17UN/rIJ7chrXU7V
4D/gJ6v3c09LLZd0YW+pmOxNXcs3yyhqvvbIW39A66PYreZ+yzG3JPds6XdRKCW0YG6jg9Tne+Xk
exqyy4m38H8aooOOOz0SqAOXCkp03CsZ/pXfr0uWh/LwG4BJfd+QWF5vP3qxmpDq2Py9q2+tZfDG
ygHdY3NJFd5qKQvATHgZRL3Scq2hpauy0bmTU+7FAIcEAIxmDLAW4tCVK9QLBayVAsLBMVEDi4JC
zsLM15+vM8OSkBnTkcV5UCLQuPo6Z09J9IFKcsHjZFFRCHq/FvZLmtVDVYGCdpbjdQBkjc4F4vPH
UTUuMxzx/t8UNmW98ebrfTSaVI5pE4fQGhitt2kwn5JFyB4aq6d9DgLCMBV6vsbaYFURTZiXR/yw
M9Zyn7LIjoNy6A1ga31FnXudRR8RPNYTv+u6MNjwgZVt1n0aJcYTaz02FavipEOi0HbMyMtL4ob4
DfJTfE0yAShE8AhTbiq0BWNAfLy3x7XXFsKgxO5ILtCg3f+lQglcDapA3Op/FgK+NwQMQkhHTshx
l7Y+0eUyZCa12tg/kPQ5dRLracoRtt5Ih92BBhxp35zCiSnViuWtu1WsAaiKOSQu4r2Efz0ZeBe8
rIaRwyOlufe0o5O3qpPNCSVY9eVg3DzHCPAR+Kqqoojudk7ZSp93RuKDU94QWOQPDMWOP3HvIDp2
YggraMfiXMpMT08tC83DZ1XPhNPEjCZAKFnxDeAluVYQBltVEpcUjAxiD0wml1QZTTSSaHzxXnM+
oXdElf9aiu86wTbzqR8w+77Box51BcOhJr9X72PQJKIskYuqdTOAtxbAhtMgTuH6ImY99SN9uK6V
V6mY12gepKd6F9LyeKTEAuB2K8cuoyP38/0NPy+g86Hp5kcbrosIyevVR8jxWZ/nKTvp5QYWTD6I
V5ZlxL4jygd4tgtLgKEC7gqXVQbLPlZRNCnQraPJ1esAbgXgabRuajAb5pM6ZGK/y3PKjsUHHnX6
4YCli2TVGJSGh+8UIUzIRi22euIdorihh2kWtGOqJRn9gMv5GElHwEvVmEXXlJgZz4HF7aQ4FcP3
wCWa10H90//yofZXSwfBZ/fGx867sW+W7qUNROpJl93fZi/sxGQtUtNeI5EGoAkJJhE22lKaYJ5v
Ayl4GzBwP/iZUc0AhKRJHrU7/dFODzIyYzJE/9rtgte5NnulkFzEgHSmWWB9pRUTk9LvO22UtWxA
Wmgie4JC6cjqbmPe+JHaptnrLsQgma/OPvpwIUQlMznb0VeDLZOo4gY5aGzG16217dhq6eWbkpbh
GyocccWxCm2mLdV25FAtY0rHZi2QsUBQUL1TqWh+Cz+ZUDUA12Txr1HciRA+nGRBzctYEnU2camL
pPcDooIvB0lbtVhuEenSODSDMai+4Yz9CJp4MLD0Tl9zaT1pwgXIMUGZucKDZJmgDYex60pli89L
3dac8jriYOKnaFg49cOXx7FeFePejx3pzAkRWudmWSJLmhhLJVLzl/DUZktG+gkKOTZfISdBB7Im
I58SRM64jLKtC14EnPnY483sLLeNSrFXRPyiMubgJkOoS3nPgiZT3kq66f/pnwjw4leKQOTI7AMg
zUYRKwyccWBmcrbwhzN2Z19POQa/k3afFB1faobLaK1k1RzjnYsBV51ADKK/VUmG2ROYOxL9oaWH
1jzuK/3GMGmGJOXC0vvy4gJO0zsk6il5SVgNUxCWjqCeP9RyvMBiquMEM/DPWugnrdm4JZYsTSlB
9M1/OMMKDjbWgELuciaXgYwjqLD0fHGyaXdasdoIOY4KEuqr5aYt8UfCv2T2Fty6dmLDe+/YSUOg
xv7OaXrKwgxAPqOprVch5k7qo54s3zSuWtbiQYEX2SiZF8Qr2a7ofyytyagQClxS38y6nKq44UzP
Rw7tkZECbAu+HKKxIKSm8cLyrQDHMiC1Tt7UiQQxuy3IMMaiBis8oOp1iWw7SR7jfFWcAVYiLEj5
d/34IoXuNjgK8o45sS4sf4W6sVwmi5Ry1mHukFWwS4PFBzbsaHpNSk/BgFIsbV7Fi7shGBviVbiT
bHRRK0k0iPzhxgzq1FH5+Y/MM4VsutKnwUGLmYggg1AUMrqlHrbExcdDumN/vm95zrkmxHYR9rut
yS5bMa7ElJGx28Q7t335c7TL/CKGii3RLmYm7j0L8/IBPTdAWuqtvE9jBcHhQKgWciE2/ADHhe3/
xqGSjP0zPs+TGKUl8djR+D/Kf5x/uPeToJfxvpFiiTL87vvJ2qbCGfearf1rtS0sRXZKZZnWg4VE
snApSHa7LWpBeDXYnkkUqY/PWVd4FsiUHGm7Q7WLQ8JaHeXguFYFcE3E4qa8WvOdrdzHnCavW6hU
SAovc4FjFsidw+saNaKvsq5EERSSlxhgLiewQ//pEcVaX3gtV76jLe8O1KTfDEr452UAgjZeZtu9
eTt7AWZFtp7cb3wAQsRj4AKvQ3OXfKux86Tz3Y7269NgY4TvxXgy0iD48w7JnaNhGHPecJy2svoC
tLozm2z9WPInB6f+PvIrzTWNss45aP/49SX1NHkk3SeegnP/bygpDq8SeS80Z1SoAwjiTRAmvYlQ
ZcW7WLTvl9HK3K6SG/myvvRWjKIh1TQaG9a+DI/tbOM08FrFTVqjbXlwSbsv2fMNcNCwXcZP7P6Z
vNB0H+jbpwd/ocvzZaMQbGaGFSDtbl4wkYVd613RC3Q+Aj2PBOqS9RT3ZfC28vwIrNnXzOH96igo
h//bZKQr/ERzD9yO+KQeb+/v5f7EakYL4ltgPK6fo3Bs/Fvw4sZx+fFH8wjKKT+oVZGsxTKdj7ly
SAzVMSrhPBrIoqC/NMJQvxpgNq6+UDozrownOZXSgNx2f3pBbol+GKKf5gavuF/i91rBy5xvpE1q
pfQc1FLRjbNObABCKiHnIN3mK9qEzSviuaoHoUjjJ3kfzNupS+W6y6MufCvjb9MEgWvH57rtDaVT
Ak2Fadh23A1uVoEK2kLF+xpGK9ASwG7501MkR8SsOdj/DaC/0PGPVzup/r37mNkA0zgrFg3BkttW
7tXokGomjbT4Zsarh3h9uNUKinctltEDmOS1bR7T3MutAlNwwFCxzIPFLwTUAusQCDdkcq2XEBP6
69giajjeA8nRGlahLFrUVeLXSBOvLPCGdcnC1DWRkadyYDzOhr5HoYV4fS3z40s5znk324kO4CVM
HfyfubqpW03cKUh6oiROe7epmCBRVv8Alq0pQTIIFypNFPVj1Y6laHHryhX/V5zO61AYu/3HW8+R
/xgV0Ufcr9a/bZ+ZdbRjJ9qBe4/9mYd+brJLSRRGXIkUo5ZQRLBH+cMPNa5ZDDIkZnRZIWDkX/K1
2QF6h1zuOAOsHh8eG9otH4Mz7X+7TBdn31srTnGSDWD1MWhOixxWL5DJsyiXGRH1ooSoLMtCJOcx
D3y1o2LcGxlTqPSTnwnp+gj5zqw3SgBAsgO1+jUr8hZmDHJXmZ+80kRJrXwYRQXYrCbLAQCry6Fn
6YQKnuHXpdKY/jNyu4K+aQwqafIJYMhLfNvOXSjnOMKSaHzmkNomDhpvaZtGZ6wA0sfNwuswTeUG
7dWKkvu6TXgdDPQB6RnLjtg+If3f3Udaw4TNXAmt0PTBzPXKcV6BNHK2uMYNYO2Kc2VqQaoZOYVz
zOEPJeQIMNMdSBQwVoRHvu5FoVHqn449y1MmX5EhaUBpCagXgTKAyhsUZP7tZylBAIobLrpSOXOb
AaY82T6tODQHLcItHQq2E1yQCXOIGj1Z/JuBXC3oSvuUEnN+3SxBoBBgbFeWqwalkJz2HMfLyhfn
ghwW7U2gvUJewMjB94qtREqYDeBwfPExJa2S1kfmBziCqx2hzAya75VhLwdsd/CtmQpTYL5mpx2J
sAz/0XDTnu1rnXIrKXWtVyrdqewccxtsZt+boJ5KGV//lMMQWrHqJc6Br9lODnXc3vXuQzsBJtmR
sBD/SnLXjPnwwvgxB2f9+eRa6y0Khd7ttHEOYbA6oVv1g6MyswKGz02fiWgyygvKJ11KrUF2/3IO
4R2xg5sKd7Bi1xoxKrMBWmIeQoYH6fQm3RfYn2KaP/ayGEAcybIgXTHylKbPK965MBjtECX0TS13
GXyMBkukH/xsUNmgK4uH2J5HBB0JLte/ASwrAh83hy8/SAeGxHPlmN4ytQ1Aw+z2hHGy/thv4TJ4
Xckhagqz2+DGLWOFLeUeeKwZNUrfuL9nyFpFC6QmqtHmPhFOxP9sYV0XXc6BjAHLsbeNN0Pdgv6J
TAB7wU8rceBxwbs1LwifWUcgyWm9Rtl0+IznkOae44xl6ohZ/U6PcR6hru479a2x/NSxgVRiPB0C
p3Xfe/OdF51R18nDrgLyjQWtNGMZzUyZAAa7DOrH3ZWGOC+KG5+dTjL4zJlSQVENAugrRbF1n+a/
Q47MKNM9eQUk2/dloRq+EPFp6clp1uiU70GObB+KXJ9xNWBjLoDKnECIOsccFK7ozdM/oh49hSs5
xNurdHyr3lD8x/DXscQtPB7S6r8dLtUw5RWide7pytTQCA8DYmyxgpluJEbu3mtZ71J4pZ1rf/fk
UykPemfyVelGaQgrQowRlYTndJIRWL9HU8ubPLF+X7QnYlDI8o/v6tlEPoAIv9Ml1Ze2Y70P48xH
OfPlnWeeWcXN+WqLBr5KTICJvum54Q2Mf5PaW3rzVH90Q/TDCeS4w16Z+NOLQXtBbVt8BduWcsMS
MPV6isdJYUGbyEX/Ge03d2/ls8XB4MOHKbFAcoVfvGqEwuKP3TRQ1oDnGDuqitBGgR9b3gYJtVVx
MDjB9gu+TrbIFSjNsmwUKWCBbTPUWM6J0I2oWrU85iLt+PGkkuAHdpaiYWR9OguFyWu2n7jd5eiU
pKZ0e9zHkBtPmTrQPoVP/vFIjcFLt1KwC0oMv9Va7raagwTSetKzqv7fwv+/rCWVDUERIYfNzB9l
FrLKeOhuZGlWIQ6ejmT0Jqyj67caqepB1q4xJbn4Rz6C0Z3QABCPp2gpXTtuHJ8l1V1dTXpIKikx
hsqaoEUOa2Z1wSKBL9Sxr4lhBco/Lhx0z96kmSUzOSU77MQme4QNhg1rwrNoovWy4EIlQvrYKc0f
ewNUNVttspq4L1X3TYmVrSc0K7rUj0X8HLfcVBFkJbE9AqHZWlg2TMuZLmIrLVAUgqnFCZ200/by
bvnxZKanZ5gt+UL7vHtJ+tWnsezcvG55aTRriJp5OKHpcwpsLN1xCq5dooH1y44JEoX/sU+sjkXK
RsUavF2/+5XRyXdwBsvsYyENseLKwxfyeeklXGy8MKC5tnFFDoYvr9ZgZ1qVbUIRy8LkkXO3Rkcm
fim1ZYi0/HTO865JdvSZf4vAoCVSEFeEdH5wPQaX/mIcaMpBu4g2M33SViV6KZ+XVucYSr5cJcvW
oTv+XGfWwYOlDYy1eOwbTf0DP1UbdOSvbpmpXF5VaB4MOmi/Tg+hVwnPmD1osCO5Zo5t/sHne7MM
eM12t1mTLqsngYLNs0S7l49Z/ExIKt+8qcOH17M5XP8/0VaF0kCbJAkeN7H8CTZi2qPWapZXekZm
iD3dPhr+jz8O3kai7qtm/hyaIidBne5FaEAwHyVgw7paqBzm+h8KikmpB812hEw9QtynOXz4zd9K
tPGrkqZJT5oPC/33nu5MIRon6XHeE9OhaFxb/RfmNtKaaKTQzqqPfWi785godSrpGSNiz9DIg5C0
xct7XdLZV3FHIYqN4qpSPjxl6uhapa0yuJJ4W/YFKeEhRbUjnHojGnyX6DakX16slWilyypikL3M
Xyxri79O7sdztWMhQ05uj2ht7Q/kPANQq3nCBt677dX2iwc5KA8OmuiBh+tnn/q4DhTSfRQh71Ae
Zxr/47aeOw96PDuSP9QsTOyKEUmUSepI6QTOarcupCleXnN9gKaKCI/ya4tGOGTJPqywxhw0l2e4
Ba3YXAkf2wuKwi5tvsOYIEi/r/7XEki+dXvtDZfYqK0hAyRPNb/hbYg167wNgVN3Pa6dE18CpSte
rWsQAJyXwo88YDQmrqTvM+JK7W8O3LCbzRYguRBzcLb1yOr0EDsKqVytoT/a5Dajz19RsLI9HDy0
JiaZIpRZrJwmqCo8beMPvEldtejAvbq9HS5lrDZ1JL+6ZKYXwCGphQok4IhTWin5MD6So41UWIm7
bLrLiRxkCRL+EgulvMhB1t+qDSuFuvS+y9CVcOFWXoPmDwGh9tXv7TK5l2H6OIQWGgi6Kj5zZ5IH
LBLYIXK0RjkKltgrQLuQ8qCR4Zom34EN8RXUOeIRwugUf0al0wPE8xpD49TRIw6QcJBWI8dIARN6
r5R6fHjhxvgKJ09uWRZkppM663Pz2F6nbNb6WiRKNK/nlLYVCZpIPduIUKH+VV6h2nGnX7sjYA4y
MbB+uZYPEcKFsBnG+PJpCnYqC1zyLoEdPjJg7Zn0Z33bBJlzZpYMuylTSZKQ916gBvCw9OIHfP8w
vFuXHoSfw6oXS3VwqnYzw7xLBOsz/dUZTTAivj4BTGe1HNdLIrltU+Ie6R/4UwFGVEfUZbdy5BPn
s2LuDYyz7asGGUg9YFWfBsc/IH1RBSgPN2D9XJMUie94cbVl8IN6NQEiSVXz1rTONdpJkMHBzxnQ
WC2rHjjxVo6POQdgRTKLTBd/R2Oml19Ma/YewKXWuFg2VdSb0bho8ajxCoQXJUARnX9i/5J8uj9K
4aNLfHwmhCVohO60TRvdRkIFvT8V3xcxZL7uL0Af8aifnz4pFW4a765y7RmthyxSPMcu1Y9s7GJZ
6pPTQ9gDTIzIf1TZ9TiHtwe+XkQc/o9YGTxkzS1IrtJcn7BQbD3wqzeygeOLq5qWVzTmezmiPv3P
Vbv3xg0MUETvQLZXoWR0aiAmpmtu9HLqfQtla+edlnAw6gfGM4bzOiWRewGwQYzQbmLL5EPFJPAn
LXGoMmlG7MvWfwRPo49YVWYOFz8DJn1ZfErVSxJKZeRtoMRjTfSkb7/ksIy5Y8DT/tthYPM8SPGy
etTSaKFx8iBs8OcUqO9tT8Blw7nkxgbR/GROUrNranh8KLI+bae1jO+FfgYmoqCPFMFPsRZQojrX
nVk8PkyBxYY8GB1DXsHCP1TQtKb8nMcQp/IQuvY1sLmQzzVHWLsZLcahdgKiyM+gkOZdWLO+O8/2
hUUXyguehaXLGsulc434QOlyojkKLaDDhMhfhjqm7XPIaFrnzKjvLB09uvhtAaP8iyVIb7esNNbz
6Rlxerd/ZQKCm8pJWoJA62sdnBIacogujb7LmTHKpQM/wlfBtoqHHRyteen3XahgUxPcYbhARhem
1lhxFICbzsn5tP/hC3hG4Ezm5v5ZzANYjXTMaf+QpeMdKa+APnHbFy80XpZZ6/G9uYdkgOFKYKJz
pCNSz71yAxsoetrdRWespM/ExInMtXjx76K5uHy/Mue3m52y3VjhWcjJfiAbFAq9OykPWN4YDql9
wdMY0X60p4nCFWigBdKY7CXdEm6ZMu5lolRIxX5mmE/r6IhbtlYq+8ociLYLY4SVIp38pquhCcM/
Qj0zYi1AgKigCVpIfVpeml4ePZZWdsdwfNPBf0zPhi7zypHLhwtSDbT6e1HGgvrPuL+5uW8wNxLn
GhIDxbglq8yxflYO1jMIJl7g2juzVbD/lvknhqxiYDPmgkYoReocU3ysYxHNuDUSpZO/DEYmoxng
73vyob7uPYopcZjogeUjXST1oQ5P2dSpT7PhfqT3adkqFZBczrzLa2qZLHAt0GWvMRk0aD3VZyBe
WkKR8nq/wzS13kUndr3x8g9Vo44bXWnRDzuc/HEFuh3kkjDte2bMyfgGc0uy6fIc9PHVkiN4KIOL
IgILVsSoK9moef/Dc6jhom7uRCjmSOz2jFEzbYP5AcHxXql+qwdYrLhrPeiaz4XC7+TJZ1IJQ6eR
eSdmX9XNnFS/gyrGIk/LPYs9P8dwwDypajFi1NjIl9+wkV6v1IBeZ2A/vgFWj3e7KOr7+0jdHZ4K
TtcWFfunn4FHO+kgzFPcI14C/biavuduGnhLUOqhBuyttWwb2hKiphhwvTXy+EysYnwFvrxKLK8l
oPk+3d3Xlz+kwhxx8DrVOqhURjHGwjh5BrBi5kAaDbB7JzDp6jvYnty0b47pGlHgktSS3/NGV5I4
JvFVbWvV7WvjHSjbguWfp6iesCLkCA1aiMi3s1WYrHJnPjBw3VPXegGAisTP4RWh52HEnRcKHPSX
8zZwuvPch68vlJZSGViJku7vYG4MG83jyK3MaoxCrMCIRQRbPhTkqIO7Nq1M+fEtojp5lH5tSOGC
G7ysq6QFWBB7B92AQDgVceVAYSLUxSS3LKsalg0kB7d1wbYd6cVsne4L8MiFLycVyLnpNW9/TudM
ONI19ry8uV4K0nbhSy5dmJhIXGr2FDa0fDfyjYg43HZ3lsNmaW7JPwTJgZSkyWN9syZYxO0Dyhgb
V91RJTI7Pstnnkd2rEy9PFkDVhtpeqULpmXwjYtxoevaSc4xTM3rN16kGF1pj9Pc2gijxs3MbPXV
tV+iHAqw/FaPziCAe5YYuAUVww4FxGiQ6Q/L49vZuXVhgofagcP+KxXOvf4BLHweZcyVPodNRiK7
l1KwaEZ5XRMHrN5EBMNd70256FfGn7/ZLhzEuhcPNJ8nISM6UxKlSHiHWg1T++kkjCyuuSdNetHr
g5TGtO6hAAQcaz0baJjUnV7G1Pb/eMIH0vneGhSaLHsI4pmcRPN5AxwT8/He33/0auz8ZF/2XlHy
LQhnwBfhs90JL9zOG3x1DYzWSR2gnKDVARHrnCA46CZIUdd47Dhear02OsWUYLJo1GbW/IfT+9NN
k/X0EiBjwwo04twJ0TcTZJoRIaNfb9D9Se3SsMPnAlbGPTzihKjKgIDolZTbnyoyi+owJZyko22H
ulP8HVVu8mvOaf5zYHv2RGoR1ou8vK3mZyJ1wNMBjqSmJmj+RNzljIB2Hce/cAAYo8a1/TYR5Oxk
x2Che5t/7aMpcU3342qbeicPCg1pTXXLLo0z2FeT5A7TODVKL3yywEbsXbkSpjlCpM7oC52yG5Az
SgUnwUWHGc/+xGRYJZBUJa8bUq4ob6vpoDV//wYSF4AebAWPCBtOhPYe8WAwCP/zAhqkzZMkrde7
kVl8i6CfzbT8YkKXKJyTUOZPaJ/CHWDsQanZjkaoF+84/rey4swu92Op72FJYbsKTrxdVv1Mx2hD
YEjt5NoSblHxRXqNQLOZEAXNOnx3k6uuep04dVil+xBd7wYxM8aqXds0xS6AqRDhH+G3bySU8TVc
VFFgLnMCHYQnoOtATzyNiwKJeUV37QPTrpfxiPK+ThxRdQEZ4n6S0hwDqee6zNj9NfOi76EcTsjB
CXXXx8iZ21VYfM36w9KQunB9g3cziEWSzAVIOUQgpYzbKPVHhWGgA4+Eno/OOMYLHcn+wGn7iYql
uSVMyyw8AeUbXHydnpdDaYXtb+s+7y0ggUp93Q90r4ON3POAT+j3MKyOWvydR9fnBcGA4Y8a4AoH
LOKvgONGhlRVNOPHxlEzPQrg2BxLiD0CPWla+H1cMQaJRRd0ZRzKgrHXCEiLBIAEY4gCCCI0jD4R
ORm30CxqdwN71egNWHrblbc766HTWWjMInKn0E+C/4apGt+mSZXCK1uicNPrIcq4GWCgEvpz8ALH
OEXipLCR45b6rOnXHeSYkiOHAIGMVfAlJ4+tdtm15URT1bR596CM5uZbu60jrciy9GzMN8QMFmS0
cMEhIdf3tKs9IAq/RnWjoUJlD74NF7iClAc1GamnBz1BAkvGbPibwnJbzXr44g+QiY7p1C1sAYer
7gNYAsP2XIffRv0+22YNuG3zaL1XcTC8mv7zm9TiQjQnvsm0l/QhM5yEhI/n4aw7La3mYkDMutzU
kty/SfGTtBqtpLJzK0xObSmIpr362p33S2BcXA4TfJPuDjDGvww4MHAk+koekal86zR6k1EuLIZd
aWwyECt8wQJn+RZXATWiQBuf7iezoCyOsZKHDGclH287eLn1eO6RIBUhLSl8wY3ZCtmyNSJ0KeT6
Xw8kuQ/2X/42vgnfZT5JlX1Jd62fERl9ogjRNVh3N5oK+Zf2oKRXsdr2mHSZitYmZsrLyIK3WmbJ
BmV5ktmhB86MoUZJSZTJdG2hEtRfN1m208b/rIU1UMe/ljJX0LG5n2EsJAF0nzrm02tyjjITvndK
ouC+kbWxsQ+K0RAGKffk4NFiKeFb/kfNT57KCt1o4rexl6vf5+N30WBDvtAc1qgVY6MJaDKjk7aC
2ZBEqBGgr+9+g/+gbO10gZPMfjsBPAnCYnoJM38mhbl7yF5mnWAzk+Bnr5AqiB5nRh5sN0uoUa3z
gP4Gb3xGBUpITyihfQoJYNSwde0Slfskx9mGGPu07WtwV0/RUhw/x8nnQsYQpxJYzBNa2Li/kne5
Wdxok49eKyyujwI44fHo/R2q2iUtTR/MHLVcbkDTZwLfk0ARxee8HQsmFjyviUmf1/2Mj64gebnn
MVJCPz4tmTjfkxKM/sH+zkvpahp2bO37UAzKSo9W930UT+btHTg90h1zO1U640dggamAWx+M+9UX
mRUrISmZmcmmRj+pjSsTwxeZsjty/SJRq+WhsSHulezhXRV6fXM3G0ByqkLOhWlznY/Ze4qHiQGP
B72DuAOw4wmjjCjZUcPVWP3Y65onvBntMMuOFvzbkOftzdBN0RZGNz+M5V3Mhrb043gxhJxJ11Ll
25+Be0EPDrQrhoXNwnhybENuvQTsBSUQaM+mbNqpRar1fQXZ82dLaVEfQdTYNJB8pMAO9Y0itPRU
sEr2c3Uj4phcNLMPN3aZKClN8exBybPoF6fgvDrOl0elb2i+SGJ+XJjjDXHjLtFkVNDzYswRPG12
Qn0ad/BvinpMsniph4KV9GsJqMPUUR5qB5kFNbf4g7NJYJgAM4ySRsHhFz6lTEBv2xdse4g+yhK8
cdappLJibJdMqwLuULSc3WYdVVYX5c0I7z84srg/CzAfFPOg7UWDSmx+zor4ChLUpiR2/b5/23b7
0QVkT2lXwnlDBh4k2L+QwTIYKjlve8241KktvRBa4NcMhFK4prR6q9tbSR0iEzUZlBbod8AUUNla
uemI2LykuT5nNrzISt4B3L5wQJgKeCnuv/5nM6jxTuExVagEMjl0DdsLBuFcJ6xjUJdpFo1VQFNY
0F+EkI4cj+WyRozp3uNBqT8P0ezJn2XeLlsirTkEn7TO1lOarPw40xkL4MG2wKyZez4fNPe7hUnG
K8wlO4a+DsPVhyxoNvJjaFBkmjrvEC0kCjMgB7GJeIL/9gXtlCbGMz/+EMGoOsBGfdTAx3cNIQRP
5mh/QtdZu9ij1N3J6aY+58cCGitB8nmfX+R5gUTIF7X13Tee97ZU0/ncrDjDUcBY//uriG9qGqt6
DfmvTnaLlntM8Xrw1NGeoSVzQSCiPslN2R/VwN6frcW4OyjZk5E/XDmlDJvyBwMjj1nLOgwp6YRh
8dhfxbd6OMUTpeSeR4cOD8Depd4L02Z70gv6M/Mkq+jkdP27klh/vHL9WAv4NfXfVU8l8fcJ1xv7
+cUszWvXA0tauYQhZ5Shx8Y7iSm1PwjZz77RH0aNTx40joHvIpDohoNQOXosJmYLfx9vimJz98IG
MZbOd4i1hEZhA7YSgmL8wb0nIcfBQbupCGqeyYmBmh/DiWqSGVRy2c7NyqTgRpQ8DoNotzqGrZSh
4Wz08wIFuBxNSc9USO6mulcWIpFTURatXVNoSq2ptXV767npi+uFSnzpxaeYq9QwWZny2cL6mm2d
0fi0QtKL4iri9CXvZ0HwwDlMS9hb3Ao8WKwOatatCgsuBsGk6ksE1Ff5UjkRfYfpOFoH5Ou/Tdb8
JBV0eUYoCTJxnuI+jdop0UN6C9USMcZ8U88HZvIvjWqjH6NXHabnm9M7gOgs/Epqhi8izncA/Rnb
J6d3LL4Y+Nf4CDnT5e5UXVQpxOYZt8g9OruoSmoXnKPscrPVCOZsxhPSWpTUL1qmED1XIhIGB1Fw
cl8sYyOriky9GMtIuaArrr+oxaG2sM//iwSG4pAgAMO1IULAW1HQrBut5SBMDKo+R22XTUL+BrLQ
evgHCXvIFuYWds3ohJtuKTKlY7tBVHhW3CVBn9oBP9ThYtT9NtfXAKfrk2mF2SDtOK2ILLQY6EDO
wq6XINL2oUoWHhuP+Z1xNEJcjD5LbHWVfF/8sqzYkAhpYPdCypfIFO4Z4dkL6OXPayt57BSjkQb4
/VC4QR9UT0D8tQJqNYbtSpf/oJQzjRWKX8HhP+cxpDJrfGoBuRoxUlzY5Hx7PddJMq/s6foQ+iff
qtGiKjPbMgEhbW89JUo/qASatM1KeNW1kXY1BXl0cOxFV/K77q3Z2c7LQIC9ByRbNyg2PrR6M/lg
kHHdMuF/HiNsssaHc4NlKK4ERf/mUBSv981FbRAGwa2XRVjiIXVDY30nBICa+fFuuuWD1sf8OoU2
CR6rvbUKCs35INfDnvMhmRHE5FOyE15+KmG5qgGgFY82Zm0KvdBBA5J3M0aL4PQgBbb6mI49EBZb
UGdjBYwxlP1APghASSMxIf/g/09mfD+cxhEld2WwirUbZb531u0O2S/QV2BLDRpaWslhpbTrA+SK
PXsNa8mQDCV4hGZoGnhFv7Xt/LPDO/W4jbnaUdTInjHiLxmd4dy/zZIEr/NtpmUo0ZFsYRpvYFt9
ZL7EdDPexOS+cK2iY+EUx1B27qrtlWI6m3W2zEee/3k3tjd2z/E8nnKs66A/OuVBnxepyj+PVKcL
jY5sGzsquHHa06+YhrmgQCod4jN3w3mkvg8DDw8yhsYx4Xti8wvyAp4erlLSGtjoBSFio30kZdxU
52b+JGuIlO5dRTEKHrU8n/9nGdY5VDFnO2XrdD4dy7XwCFpl40riojoJwwb/XhdVMGI0sh9H/2l9
VjaFuhvAUeKrXQd1/21Eyw0+dup+jzSVCZBd7zFDRbOoDtzG9tup4mt4PUnaPxtpTLa/DMUdPfqK
ntUntTFJWnWHB6W1V8oz+gqsMRUqhjCt17NzmDL1FHL2VPscRMKkgoFZ7JxBauLuSg9zzebC3r3U
1TNceLvmH4H5IrqleF+n+1SBZR2IfKbEFkY1ORjVCxCvcJC9jXaKd2FxOyWXknbuzjfOfdJ0Epzr
lxmDe5nyORr1p+fqLsSs3q+xdIBWOh280RfOU/jmGhRnbKlsqDP6+Jz/HTpPrzeJ7POAxzuHfBPy
0+MiURgMg/hyVQVwMrGyeFhbLNAlMCYSGuyjYx/cEevTCsl/8htZ4AQGk7TE2HU4DWLmIxzmrN5i
Teg4kfZCpC+eaUTkjSgd9ToYvO9wJuq5eGg2kTo6mFE7DWgUg493ChxkjkpVeiumB6QfpGJYqSnk
EroiqmTsCo3MldWqmfy5bDXzXgmD1jaVaVa/ahqSp4DANS/Lj6qDEcW2L3Sdp3RFGQNcfCv3sopH
dvGuK39jpGqtBOZSNJMz2s2gwW4Iar0FKe+xGvfsjkI+qGM5lIJUUMeXvaIgJmyTqz2IhNOxZ/kX
VuY6CIEZ/Lx0It40kHE8Oju83M95JAgNvDj9D42uub5JD0BqoqZ7hk+312caoZzCeLnEZ4Gg0YJQ
fuKeCb3LRA5huHc39PN470IMcdXXTRY/7F/V/E5VtRZpvBA8uM+Scgp0YesKEewp4zaN6G0U2zXA
D4UxRyjl4ZM317ZXuO52Ig7jDh95msXSBGhiWnAhrAwghjpKASHKMHa+PfYEGg/kdXbdMbHEqKKh
CI3tKaqerWwDhinz/qiqK3rlPdjweF7LfVqWAqOM53HqSYJXJdUSZmcZo8G/RveltDv5gDFl79It
sgSL9coXBXrm+6PUfYSWTuxIuyfT3nB7lqCycO0C3g5ofl4Cu0RAlxaUtNzWWt9FmDaW01i1i44z
pkWKdztdl6iOccQv5zm9wC0sHI7HyjyjA9OJoI7JwVErp8DelXSl4Rdznm5yehVmJT+qWzOlQKCh
s3EXWs2eCrUNYpF4hSjnClCCXyqP4C6Ik761diCOLBhiqv0B2GzeDCXRoDdo9iVxlW2hQorequ9w
dA8fVFch3ehVrmBVsGhvmHKE+sSCa7UpwUWZ4yiPimaDDcXJ788TyEK2+2HFdCknbleZKoQdNUSO
v++861lvt75oM3c/Pvuk4hlv4TPkTrqtDvtqVA9PbcVIfV17SLmid6AqquR7xJ+sFEfMhnbpoQtd
TUTY5Hnu5JzvT1P0K+IF3XDaUyCJpArW42yNwx1c6aZ3g8lqysoyjYOle4ipT+W2sGdq9PRrhC0t
R4vpaB+fYKEez4wtV1YSGe/5D92eUWNV4aLDu/RgNh5tSg/Sh6pT4eZtz/H3C+4cmJYT16cAcIwZ
xfjBpyCwkTzDzMIPxnO8XQwhgJM9lz5d71unDrZlpTEViWdTKm9DXjRxuqQfMzCagcYYQi9wUj4X
F+eWP0N0HeYD/wxP/db5t0bUgNm/rwR3E12jGdMAQI8uTCAfk1w4u9xN1Nh/5Qf/xmBGHMJX8tts
HSSlt/WDUNvUayuLe6arD3f4qCb2j5Ue8x0Wv4F0zsggFE1FH1zJl82QHSjZtlwCpObuSR0O9wQF
YRwT0rDrje9fSGiovW37sociH2KBNLXlaTYImav5A6RmIdBbDx053UCCWE1Lfz/VO/RRa4JcxDPW
SiYRKjbM1QZrHyZdPex6vysIB9wNEaIRH474WdbPCUczDAHk50iPnzUz+UyL7oaBkNQUH9cwydLX
c8mW2nip7AedUdzRv4u5uOL379IQhMN3OLhO+ND66LVUuh8Y6hJ69FJ7gP5ZCXiSZe9QBxJ5fV/J
Oed1bsggx6IqVnD+gP6vdiQGwzmz2ZiYBdCMI00k+xLBuDr7b3mWqP6Cjrk0UvkS4rFju3Emttp4
DhStPd34CZjnpJHB/2TsjGcO5R1Mj/mn2I4f6eR9pfU0fzf0y+UHW+XOklRiwLdf1W7iHc5Iy1wJ
LgqkTBao/jjcSXPY3BbEZQiwkusxbF+bKE0QwIo4O9eCTWbuycCCxj33Kc2RggNgv8Z13pN/tX5X
I21FSPnNzdZYy5p4b7jSrQHZzQ9oIZAWpvdwp4qjUaXn5wp16hY17CEO0cECS+LMLVJu1Yy8vt5R
qMWsIoVMuncSq99MACe02t1Ms8MpsSxdN558MLbVpCvS5xf/UoaEy1G8/RaPhUIs9fehuKzjG7c6
bjp1f2bOLp6jjVBlfuaIjJRskgUTQSVkIVoNCH8qsASutpH9nxoT/ZwqH8at4IU/Y6DKy+O/Sern
WKxK27MMoUn2oHNIYWgM1cKKbjyNfognlXIvkLkn2warGhIwP8UNuwqU1wdHolRr/dXHOK3qqZD/
xlKFplPATLocZfTutXHM6CB0mG+fza7i58v+YjGtXRRTb6nPDwKImUoLEo/ePOikW6XBUMLpjwYA
gXO7Z8UZvnUwwwmmUAyBhmtYgp43VUgA9R0K1J6UmLGNOki4uFhb15Z2ZBPj8Y8kiZ5Bx+06EfvW
XURVa1XLDnyAjKk7IT2PRMHbWJCa9muqOyhhGFk2uoozxhfBv3zJfnihVQ1R/1EDW9gKkaoBoz2I
I4HFpYltxVviw7eEmHWVia+KnPjr9Spw4nyYuENJ0vLG/N7Gfvaut+KVDdP+EJfki5sw9v58wkTA
Ya2A/Ykdy3VLtTWcjxOF+k7fyHvVgOtaqonFwPPSjM9r+O2mjyIRTw0S+R3uVfnYq0c9I+STeYaa
ghCEYQQrFzq2qlXNXLAMw0JXdGh4EDOl64iVF4nwP2x0abtRF+28iQOnSVxySNd1ozSbSMJwLVgn
7THMdubMiZ3Gj02lrnZmqOQunhcOlf6nmERpdmTCBo793BDlJ4TQbEAfbC73pjtyACJUi7JR2ym5
UmH+FG0oXkIKYoI4hdRvWUylgqh5IcD+JJpanqajjzjw7moqDz8ZgklXy8INWuj2LY3xHsF/IUsu
Sx7KXXmlVVseTPECk5VeANQjAA/JSPQeXkfL2vL7h/XJnJE5h2mfVIdEO0EwQ/dvFbYrZwNWbuV+
vLHkD6eu6mIJWoaqOuh8SHkGR/MNXE4hBe/y60l4tPXEMVzAEW5DT+MLL+qX7jKoHA6eC8p1EAJ5
kJI7PGijnxlxVaBn15L3nZlbPHoZgAdZ9da2iKqyS+o5wdL6UN1d7OK92Merq1pU+Cs1yVu4frPP
rFB3xavqCOqmVxwCPB+PSb8P4mPfdV81tcqdTetGq1aZXtoP5a1OuPgcx2530pfnFnS0yFF+/yQ+
0dBkj8CJ6XQgP5k3VVQn6n/QFfqZMsd7y4CXUhhNmki0bllawniMGVN3LLqWEb++BqXwdYr5EoRO
9127iMmTpGWQ3FhNWR1L9cgzm1vf4WNXVSNh9Vbb79cd6l1KY6qvXAuke5HT74vs7wha/4fRdP34
CzNSrFDZTRZxYebxWqjqrNhV5qp7VcZbNq6eSiXn4jxyjV7p/jgXYjt4RewM68JMCMZhcoRdBHHF
w4FUQeKvkZ2bA+H3DgdjHgo7LSuWc/z5Y4/fiFUH2Fqt9/oDWyyn/jhcLF0kWjcWI5NeewUZ6szK
+R9xd2oDg/SKG6FOmq2tb5Vrb2mX93zIKjXhKvHrjLofTAygCVDH0qO0tTH9h5oDRl9VgLcfQG49
zbkmFXGC/O6CR+zuuaBHfKgQWdVYM+ge/hU5oCZgewCESy+FAZ8nTq4wjJg7IcIME8RfdF9OSK0B
c64RQlRZ6kznNFjSQaoAsfZ7+/u2vrs+vLCun6kooa5Ok3wpnhqgh9EULcqS2RgSIohAsB981/57
kkHB3qMh2ZU2BwSCSBke1SIom9PvOunq4HPSNHoW4qiYQEG9joiw2C38R0i5Le/JQBZ0fHbQcRUR
VE/cQWkHf/PBGhCfccz01scujoPIvyiP5Ass8x+yIIQFpYdUVdSojLcwLsMX7PoUEzjjTP4gjkWu
2pUHnZR7fL8DRYAs8uMC4nJ+wGiUhSY794J2Umbpv7R3kPFIagK0W3H8zUm+3YAkf6c/bbOKVgL6
J5Gz4hE/AvX7peGwGStNHkVtPSPdKbdTJ3+inR7HSnzMFTVB+rfJxC0ZVmzlMztBMl3mBo3zWfr/
856OqimDR/GT9rc1AYrIatqKKY8sU/x585BLn39foJEkbNwN1DQee0GKJ9G7xFnmpGhNNaNpHm4A
+oV/9h0/rWf/WZy8k/Viw3LeqtteExBuvmNsg7NAbGc/fXTlGuyorDcWSIxjjDs39NU8Sh8OKDXr
7v+kYTVikIp6Azs84zQhohoIkycP7IOWg/OCYBQqnfpFOptxJFITxh7fG/9F8BCmAL/GxZhOb5tY
QLa2fdxg5S7+Zhg6RWf6C8fD3dV884LYBAFW5m7s16YMZx6dHZyNFhtGUrAIZOT7hDRpqvMS9fQ9
yrXTjMUQCHKNLdMgXIONvikKP+Lpmnqs+vo2ShTZ94v3TaCnO6Tk5zkZDWoYu3zRFWQHKjuN78ou
gGvF3/zVw3HFsFrC8HCcLbEeTCLhlKPGIXmfLAWlLwq6J5840zoWo2nuPfWa1p54wtc1T4ytsFYI
qVmJCRkqVKulRUbc7ZTZqx7tYt7qE32K+eP8k6YjyZrUa+uMd/k9iIh09ZU8YrAin9Rmr25+9CCP
3S366SnzrSbmJPEMMt7l/aYfVXFSON1pGdAeIr+UnFvihPR3sWQoGCN2VfrpOCioWriwHuQokHAk
b/kTdPd41caOjuP3ZcHVpX/RJFrRpvFkPcz9En7ljH8butQn814+gjgCiKoyEFlRS3y0YYkwGEB0
k7aWUPqIqiJURJXNdGxaVLDSBIvO00kjauKLs0bGXLVwrurNhYNtqYEOlpAJ+hG6CcG06cCoKjT0
iso09w0/vl8Ycni2OI20G5OMgbRhCNMsZbjpzSGQPVyZFM1PftoFmQrdfC0vHreENVdn8Wm25Q7R
d5/4gNfzU5VNVgP4zwNglU8frqA0txoz12Lkw1odHj4PMSsRT+HrsgBlEY2LOA9/7rgKedLQn4NN
/1KX+ZdEv6m4vkhJK/BHP3EtPiJYtsFnxrs+ISN8b+u22TMbMv+GaupL1RyW+QHlFY+7rdCu+Wwy
Qe7hhpuu8GAuc7HPlXAI5abDlS5TNxYpCZjnl4GEmTAHObdSFXu/eyNAPaAX5Ul0408/EnpSC3yQ
JRHv848fzPeKksym9/bX/ybW/sVity49CMrFy92kH5eBci7x4AUetSply2feO20/7qpvGab+UL1B
Ix6lZVi1HbUsQuSaSpX6uRigBXzp+6eqeJM7Gj7YJeqcDhMLY2QAy434YtQMvZu+xY+OD1ADhQpF
omDXYPcd9hdDXi4WGw5r29GlxZDTgiGk5uyOxmGUwUJ1Y4dO1r9cDeTCahRCPZrOA88xEdrYHed9
FkWzg6PzToplK0CWz/+cCt0GVp1K+xLreFGwLPl60C2Yeplv+GTU8ZwizceLX3NW29QC2dIIy5cD
iPBnki/tvtUp+cJHg3A9i031xeTf7lfTS4pzp4uTpwMNjOVzFF/t6dgVUp/vksyDDgJu3DJlzRcE
0FTe+IKRYm6to+O/jdyFvuF6tFIwFOHT5AQL/ZsRwNT56vksn9T005LYWz3LaCnWh6z/4guasAIr
V2VpkhNAD6j5b9gC8CdYdnRvcwxl0JZS4AWpB4fKpGcTk5Y8G/6+kzbxniVclEhYIWdS5rNmvCDs
Rv8S4jWis3VH9YpqaAeYmFjAQyEs+eFbS+0WIuYsWXeBQ1X1A+kRgHjBJC7SRfQTJ/df9q4A4j+e
aj55FVxGgQBRqqrEjCnbVpK0Hr2jOMsKfJ8LE4kGqgYeuwmB5hgeAmS4/NTSn17rtHdEpWdCjS/4
BJavlx6fYOLr2tyqyMwa9BUA0Gqk+JG/6uAKAPHqIG+Ybga9fDhHDBO299j8pfWw4iDyCls+hIg/
A1fn/PKHogoTDwsNyDvnpFcjyPzUmQ5LRCdUSTujVI+RPh7+CWEDrNw4wPAFuUvizVeiIc9jw7/j
JeqCrb+MCbwEA6yUqDe/x/cj+nLRwUVwjVwPU3tiFtS7h5oIStWibMk90Ier6eRIZY+l2KQYUjtF
L0UEBAie1CIgGwbJvwKkIDZreRA+OJAMt8Vpebh0OlRWPWovDYmiAHL1knW/EwRvfLifK91oH2Aw
SNTaZEZ2Vo9d1YEgEZMjdm+7MsC2XRRUtUtheb7z9npjL7I8foipYSHygmvE2Is4V8jPnfcXfR9v
Lmpp7Y6QnCEGL2c786tOCjmJjlV09H3oJ19FFvWBHnArDyypffSeg+KntIk96RZ6D6AYoSnScxQA
uWDbAvhNiRbIipGAJKuoWUSLwQBDtrGet168G+y8FHaTELWvUdK1Q2UJFHmeNrAI1vL4/DCs2IPh
HPtFVQkvfMIz8g2SqMqWjF9rPNDDTOrnh4WhqVx0Mv4JrG+bA7vCjBw688QzZjdZyhd7yj7eGJTg
osB10Ky4V1N+zKWlGyyWgeSvf7BJJ98cOfj49GKWknEIoxiCC4Z1ntZnvIsVhRTQN9xpDZlFqui8
r2BdumMOI85Z+VSQ/a3rculcY9KSdFQq+ytKnMCkF2eyzePJ5YXuaTW3kco0AopIsT05QwruY7Hw
Minhx4ENkwThV2r0CsPD1yVo5ZUaJ/XsfXPQ5D9BLD66xre4fDGSuO+J8t74acAIrMSxOG78fG+C
ldzUCxU8C73GLSPsVmpZ1Pndq6bfzo+cRjCDIJw1xCoMFXlWF777Hs+6DGcUgQkDlmahnIAR/qb0
eP2f3DTAMqaQJT3sVnDhLX6x10KKgqux9n/CsajktuH4f6QnxBFsTNce/1WtptSQimRO9UHuWeQ1
Ltv576Cuus2o67wt2t+/jsI4wPaC0VfqvoFxYZ2fFwWkk1NBL9IG3oFhQ3UN/Dq4tTA+GfZ2leX2
RA2XFsjQc2vFNVx6f3bjybKSNCgQ56JxPjsfpQhMHCdklG0wpOAqSXfyzN9o2x5mdPz8shhGO4jW
a1ysOMjkJ175882QT4AnTB25KQqZCDLJsImIcYqhU01NbFINzv+DSu5UzaVpejHSddcHuo3jkHEY
tyP80trns4HX67Pk4OY4LQoc04exuALY5ukDnwVSaUwfulsrHOnSCMACrHeKdriij0hkduTPHznL
BJm2ghT5vjSTicOF2Qpc3RUOVMairHP4tJEJtwTmjbBu+n8aoS+nfAWc2DquDN73Fuf04G9uJI/Q
Ui1ZMo6kQLiww6yLPiq/5ADIGdmnk58KdlLxc4+6d5XZ5M9BM2JlK7KB+3att28c8D4bRYpIwrTS
PXXSjTHWizpaQNMu9Erac2NE5niR7HVvBVtagnAuMKLb5Yk357u33/9xetS3fYDMd2Idpan/JFqB
yc99QD4hIZuirbC0lGaAjvhYulSrDFTf9oFwj3EjfDVo8rgJEGDWFmlWtVPdZFPncafC07oMONAr
hdIl3WG3JtwF0Ut0zv/+q4JART1wAZLsH37q0TzT5DSqSkajnYcZum7SL8pZVtXcG4hb+pXBBYvy
VrjNF6tugycSFgPF+xRfspceDcNDpT+DAqz3ybvGl6Vf9/vmD55nLQJFvSAyBmwIARGV7frcAQ+Y
WkSDEup1VhsEasqRc3kquCDOIJ0t/tcqBR1N9Ej/S+fG5z9pF/03V5oeRYqLS+e7PUsuCwDXXVqB
+zhu+VvYkS3w2ujWMX3R2cTXIaRZ18KEcjkmrjxW2MNa+E3HtxhTXXlcRhVsTposDnCmuSeE+5hU
oa/FVo0ElIQTmWDPIDcykLaIwKf4mynWYCdUvTswWmXcu5PwEdGU/Mpadjr5IBLsVJx07dRZ+ys/
Ro+bSeD44f85RLF2+4xJOsXAEbU9mmgzP288K0zw8/UGppoJ68i29y2/ljZ07g1sFrP0SXhVc94X
fgWAX8W/UqIdRdcLzD8xgaosD/DRfpR052VPBivmUGQOfbDMQWUqShOBXlmODYiw8+rsnyOa/NSN
B9gTAM2DIk5NBPjIFkT062cRPNulmqpOr5YNU7bahzDAxJC0lAPpNi1TsnLByi6P7cvbOwZoL9FE
g1eN7WhppSrvQwCUoRAABqar5HCXG1I0PldN2JLExyBLeEmYDwcXmEP1nCBCfkyjev/R7xw+fDru
Elv28jCPtiEL7LCJxRLKvhY5fyBqfxr3suJYj3iSlXcWSiXqDI+3obJWZNDqOWWvb4vx7xV6UvyQ
RdttwZk6z7WUQ0hakSQGsEOXKkDE+68yRUbG0qT2GNQyBd5Y/JmazaElRRP1z3tMnYsggJMZKubU
KNGLP2fdMeiN1Qf/URyhqlYNCoEd2Hz9upOSZG7AllHN0QjaMeC24tiJknzNUsnL5SuzVpEdq2EV
ihLJzl04cT7eGnq2tscJsrkAxIigUafl8eULO1oJJqIgjGEHgLfow6A5hFvv97zKpxjU+o0akF9X
Nscr2VN7S3YENG0AUILBPMAzJyEtqlcIE/8XcrY/MZHqXb8psFEY7j8MYMnGghSjnDE+FUFjINhC
w/OyEtWu4LeWX+9LQTG3L2tKDVQ31DLSEXzRlM5XLb3vnJTHTIoozut2GPMS/fgDgjdJ82Z8dLj+
Ai4qYPgG34eNvTrA70Wyp3kUB2BJDEm5etTid7dcyOBc9GamJx9qkc9hEzpaE6tMif2dtq8OYeL8
BzEX4ioxBx5VMMF4NZ3ejNPE807+L4iSePAWbKXMl3RircnW/EUSevMRAMql1DBOQpGr932DvBt/
wiR6jChE+bSzj1ATrhu0qkMiCb7Lc2wXL6r9raAhv+rXgVm06oJZScZ9bKraU/xvVHBu6r8t6MHu
RGRajrF6rH7hlcVmWaUd8MmhO5QYu8gUiYdDGdUal625X9rO8TxhfxZX9OGw7L/x7rJnC9i3slRF
8VoCWKxUs/K16GgmlJh8du2j3gh+tgnhPnaMruvxSIkNYhvAnyqgz1BZUWpd2JIsJXBZAsRWMgjh
T9YJvxMRiNmW+ApFZYpBJ1v82a2wNLsk9JVnwiAOhqXI/84p5qaIW9atngPar22PPsul+GLww7MD
lpOrE13EiG6nfMZZOFvo3+J+YCN8Z8jtJEOEU3CKOeBXUUx4hFe6e1J6lxsDKhJB/93uzGXo4rki
iJO9je8s6PI87Jm+zwP+fxH9xFgLlrB/blNTKtFVvSabtcvBQZykeXmPCy4VVcLzaLZqZDZlmVLW
3EKfBjssK0ZJ1TeM0jZOF+bZyKJYZ1DdLpZoTJoeMtp+EFEn7Q1ZBTh9btq51WM9qMcuS5IsrR7W
hI253fEiMGQvKfOSwj3ci8uQFy6jgCXYQ2l2HizeIV55mU8ZygxjRpv0D4I/kSt0gnPxJNB+EGtK
dJy/plCz6PVhUPM5BijnFLcC/mIaesy8L4Z5oZHEimWLNCXmJypIgHQ3LLll5TiMY71zpoweCYdH
k47HzVxjXnPgHE/CXK9iYsk7Q2nqDTD26inXFc1ZCQyn6+RBAxbIZeKCcrna5MmTl01mUy1ZPA+Q
fkBl/3ul29lWnERqWUxE9W8BAGR64c6T6AD/wwX+e09nyF6ehOZP7d/ZvQvwNs++gouTWdJYg9Cj
vUGWn4+46yiBWmKOFKIQhBS0ZEMtEtJsZJkkBAluCAzodA+JI+NF4vcCoyzZ85FJhpQwxeB+L2ge
MGvJLDgZJiF9UfggqpUkWLfi7oM2LATOugBuNhE+bFmcQ3tLPnDu9AdXvlFwFGkkfYYFu04wxSfA
/E/zALe7HXYEdiAOKInsB4Qft3G3xUvPcXk5TWMpXRqKJRHQY7xwDuN7pzvWh24XE1ZwI3FZkfGE
6I9S6q5mfwTHoDceFOqHxgb0k/ZdeOQv3eb1b2ZkSh16xCuNp5np3Ru2Nio6RG0CKSwWzwCeoUmo
TokUq+LbRa7WkOW287GvVDsISBmJ5PI8NB/2X2SYGFiy7Yrj5E+2LtQ5HLeP9VqTdG28ZvkG4LIy
IyyjJbWXJvWpkVKY3O2B6ixWQdXUZ5/aXin6qi0wRHYvpJvyYxKzDCy/2CNAB/50bOYUtlh+UTv0
MoaTvZf1H1hFWRr+APzwJpKHx+S+Q9FKFUj3nMZF5PiaArS1H5V1gqXYkogSrWUwMBr2uW8d7POG
p+qaZWepShtvVatTT6+2DR+sRKRzMC1qH5L4tmTD1IaonkyQiv/XnY1e7caYKlEKO2keh6EKZi40
pQnkJ2aA8ozsAJ0+9ZjDf6bW3+GBcntIz4XzqsZGlMhB8X8GaUyNxZ0BWOgLKifgxEA1tszg6O+i
HBDte5jjp5xLHG6fAmnOZjiXUe981jSxG1+celE9HnjwelpW+5Ik7RglmN7IcC9zcB9hCKph+eM9
vMov2om5DLYy8bOcizw5b4jrufitNiFmrVAvHsUgAJMR9nvMT0R8xG5WJxpT7ZwFwrDrmAzgkzEU
Wi/p8hok1cw7BaDdyCAmtFN8Z2Nr9PwBPrhFsumbLRzf6GX2+hofIXw66HTk4ll/gc+c8rmc0Avn
sDTDQogub6JWFX6E+lGtkDflpGOKqtARmFX65FyiOzeszm+DAJOrqP2JPQXjfnxO4obeeaEZPigz
DMd/Lsm6sjHHP3RUeyp/82VffJeI1Z8nuanqAX5dAFcIAvcu41oqMNWQ/cPYbETHZPaGlbMAe3qS
TB31a6Cujds/d6EAK/UN51ADqmUIDvdmKtPl4Akz6TpvVbB/Tdf7CMjm1ojJ/tgPZuzZssl1ze8V
pItoxe9rqfMcBd8jcawGOlN/uyhTMwKu7uJI5lzzO+xoJqCkzYo60ioadTVeMFmZxjUt19DMNDgl
dvzGuaCWd+Mdh+IAtkcjzTmL3qhZ4/Fg7Zww/5ZNIGpfSKbAYcI3TH87oSCFFTgmzlEI67BI+fgL
7DEDnAkarM8y/Od72HxJAbYkUN0/1OhgQA4pYUf0movPv+nvRAr2ZpZmf29T+ERAFeg8qoCOi3f3
ssu8Amzw2qDVHLwI2iycSwhcjZ/WIE43uXrYdY5fhCjvEb6gd2O59/TzMfPckDeBjDIVeqWUt64X
2Ycp7o0sdJzyH4l4T8uCkH/PpAPSRci6X1zCeeMIQSOrvXgOyTtN1l3deqiGgyaP4wyTtEZHA7hG
R+iWnbT5X4NovvlQASMW1Uz6hma7iCblfl+wSYZVBTVfCzfbWmq9YQTnl/gm2aJznv6cEXIKrRhQ
u3wgeuudOfzPQ0/JEPiIQCBeTUIDCKV0cuLudpJlwJGST6VJRzWKKgfn4trvThv+Nn+dZGxkgJEc
5DXjAZJJEMHA+knhO5git6BZWzgK8jMeggLb1rHmZGcaCKIWw3UO1kUuIt3ppAckmqkw7WStEJbh
D80KDfjy0ZVhhkiKdv0b2hrzSKXv6ew2iSvHbxViEh1NVxl3zegzwXSg76C0OwgXGMH2T3b0pLw+
6C5dM3VrpyAZ6I/NZFNIrBN0EPxQcqU02bLnFyYBj12ZfUDJ2RuquOvRihGmO5ynO3ard7vkIoNi
EZ8TDvxh0KcXWQ/v7/eTMLng4NjN1wh0RfjKqLwrJ64x0lKLLZ70ZmraLOynuP8p/0uwBkszWiKR
xKna1nSNMeuTYLm89z2TKGF7/SNIptdGyqRlG0FRudNkVoaetPKoiS3gK2GnQ+xp+ZMIj4amoLli
DOI6+1J3ZAwAMVn4l2Raj0tWR9IpZHO+dDUOWcWYSW9WTd4m9wqQ9x9ymhkVOFFfS1otKBFC018/
pxK2Z4pER6xHBOWkET8qqfRWwy9ZVQJFGpn8DG8m0UlhRjmoqrYtLy/4LfM4CHATa4qf3Q6aeH4R
KB7emeSFoZH6BNGyCAH4L7+dwT/bIqWwAiL8nKXOKoAssFwrg0Df7KqV8N/wYjeqcDgX3lBqjeOC
Eqm+w2YXVGilOYKWvWVnSm2E7XStAExil4lwoZsGnI7BmLdEhrf2JV3rbe8GhvEG9I/nW/1r3HxD
4uItCdcrFUu89VxmWhCLqz8ZCStu6J8f9oEJhFl+k88+tO7c7mctNNvbS4Iu45bZJCICSR+/uOfZ
3OF4pRt6IzuMnWGoKbtpMvq5nnyFpnpRXKsVsxb5qejjMaCa49wQD2lawctivwqVjj6wo2/RKTmg
ZZrldTUHa+RJ1/bW/kTSUj91rLzBtMDpMlGu9r+eRay2fRSKnDae6xPqmgCwjqHNz1yPiCfZL+fT
8UcMouViR/HguaTMa1e5INZJTg2YgdERVeh9P1vXYbdn09W2phu/N4Z4Jelt2ALgWvZKxq9i2ALv
FBHPd8pKZcp8ViA3HwJ5KqmOmW67pVhMJ6bnjgzUeZLopRXJK3u3dRyqJ+yGKpzcJmEypRF2ESH/
VEg4cpHjYcn2N33YC/1xxrJEoeWqIHA9Dgbl5t6IGzf4SkD0zUQY8W0xAGAuZhPfqdNSYmwB5qHa
5v4RJW3fP6gzrMZin39tSVyMjX2x7yad8AGZkRXzertxIR8rVv6ZdIZH7FOei615wX6B+taDhy+P
H1r/2187YYrpJ+ikKqHPkBmlj2yz2uxBD7gGMTq/gj8SLLCkfq+hnFdgSpnEEq1SZY4fFLcLndch
iPchw9f6+DxsegvhmDtW36zfwUfBInc/PyrZqv6O8SzClyU0CorYuckpRYTdS77fcWftTPvi478S
CCQEPPeEQAA5I89tsH+urq3nOL84p3M2Qqt/KVtpT7VlHOm2p+oVB1r1Y4lj9YngkiHEctW3Ba9G
zEjpT7GV4ja+9BfVzSBF9+9PPm2u2WRg4jHnCbilRFgNHE0HQnDXBUssOSUrENKnxHA4eoqxolQN
MXtJgMPKq231cUtqyiyb5slK774lID+w7exCgG+AQ/RORQaK7gWt2zWTttSdryoWPFb3lRhpVGO9
T8s7+eQeqCla/G3peFNHu3U3Cco7XyT/s9h1zrHdRznFUqN51s7b/UD4zrUax0Anf0hP43ofTWKZ
oRvpHW2Q5Oj6ne4C0oaebxHAono4ofakSy51cba9lezUzAVgn8RZwuMgVAz+BnR+pBnPkr8fX8D/
WTPribcmqeGyxd/8sBpSDjtLtxYMfoChw53pFg9tbRMQDtWEPk/V4FQKYP1e/AQwct95UaoswnkV
Mb7x14zSkT2t7sNNgN1o/XVXu6chTF9Ca+oXV9KfXCyzCcBCPVL/yFOiSIGWdZmdW2EcUQK4EHoQ
uFNfieepXbPUXRdzzYI9G/DfGWpzL196MBoOcCcdyhcRvqhyABN7HrL/AC+c90siTqiLyEnfVB6C
BROTNzFJ4g1XGr+OVvNbBKgFoUT2btM9wFWtqLja1+htEs02TxqeTphi/cpcW5Ng4spUmmHIiPef
djkJ8znN6EPTx/maNjVFZSeJuRg5/BSaLJ28z0pB7Px/t1ryKLAhAM1WpxgIwvM+vn7afWXC9fHy
Ahal2fiQNtPPOvE++I//merni9CjZlyl+po75UqSlp8CXrei0+jZWQp+/LQ5LuqmE90BOpw/+sU9
5x6OU3jPnZ1qAT12J+bSquhnU+pNUtemN79M/ZtBbGqqhb5f9DG+zeOm3iEvU9A31wJFCrtn8JPR
+SdRO+8qlus8rhikROcSaG5eAp2ASs+Ah1llVveq/cnBHT4oQEiZnfz4Skevidx+sZoJkxXZnfBs
cRuBwYMdUfoXZzK6776Q/+plPMLqpvYTt4UJZicnCq7pTCrI3TCoikysATrtRbWRkXx/YcgL19gF
kWK+Qii4s1GYsmxSR+TzywDT6KiRV8CPrRzJKJfseJ2D2oSlj/UvSwRdTSwrl4Sjoxo5x1IPZ+um
WQHukUk2uRCkk32W+X4YB6e7vASxCLtXMLz1CuYKyTvflPt9aAaz058PULwzfKSJIGR7mrMopxMM
IM82Z0lkht6doGjf8edBknWFs+BrcP0wzDjLO2k+XOVcP3sGIkm5aYd4KvNKvi7A78q8MiN68qBA
SGJjNQfr+k4UH/ARvx5zAOLEDROQaZwivYh8pNmbdALrzQ06GQ8gE6puQ3sxCyTey09vEFLG6J4W
5rF56Y1dOvFl2pK1+wyzWe7G7VyVI5mOQaMGabivVIquwhO3qwh/Uwk5cOW1rFJbukcsbjHqmFG+
PZMvXVs/67usPgqfjqRv+2VRuF5trPqm+kJG2QPeNLbM1mIuQUpSJ5cthxJVuby6Drtb1MMHD3JO
TcZ+DxL6qOXFCCTUiIgBuf9QSsiZfIHwakwZzrcXuBA1LxPLME8amJg84ZblMJSzxOM5NYULrEsO
Ml36dByqgBscmvGFFEJWfR5eTo/DFHfOziDrpckp6AfLCOCBfrZdqi54oFFaICQlt9yhFqgEq5A2
zgNLt8yDOa1bGc/Hi9pcccTCIK9QiWjuekBnl00B/bV/MVY4soiEoKb6qWUGUaqy2lK/HFNDf19d
h20N/XlflpmAKSSnsCWZ79kfAwkSXQWH5C1IYBPqOH6TekI4x1lCB2TRQZ5bO2q9wqKdgMwXLdvY
9BGJO8btlcb1vA19RLlThTcT354fngBoA2ui9kY3KoisjcmineGlmXO/sP1vX+q4sQ7VXOBEvCau
crjHgiz080IdJ6I0/hbC96Oo5/t73NO1uDfRWgaBOBMoCNnqdyJDwMpfMh+fsDdLnynmjwzR7OZN
L/MgaMQa94FAfoeon5A7KFcKCZjVvAhPPgIr2/CoDl6Dp2mo5QDitx5KtMEz+ynlhGggpCjfcQBa
TIAmQ4BaW5HvKVaeXNICSt3YsGiYp9zZF7bNBegS0P4iyqKyz+6yp+fOkx6kCoNU1Gd4+b++RxRs
BkF+kwPqGkS0mCRcUmQNkn1LMhhfDjdsDlzCkaTNTxpTYDTFOIaCKoOgeR1Ig/qQ646vMYB/ELph
BZa2Jh1oA45RrKRLeqByCZgXHwVmQ4uzgsSVBu5RraHrhZ7E9rQ/Q0Ic375NVqhDF3oLlpfj+qGE
4PBS8yng5Fgi2YnbLWlAb0RTab66UyJ+vuiSMhzq7C6226aETbMeiLcKr03e+HAC5iCCikF64wKz
jbXVOouX+MwUxFJ/loe9Wp9YmqrutnS9iG/JUuXVggs4WBasHh80u8nbYbviU+fGhl5reLACsNfV
5MzrelUgEsk+JzPokBfYzOtkA4qtfdTKlxPq+pglKolPFeL1tiQyAzJ19n7mOiGNZmhs5FqPEUQ1
+H9ee3JN1/frMBR2334n0Cg6Pot86CkFoS316Ft7SC69Ci0B704GdxweUI995jj1esp0aDRpxEoc
GogMljtBFI6W50zUVRDayUgTecpvHC2pLKTbmPPffirlbQwoATb4W/LybIJG+CJuEGVGFXmKlbG5
Gw9AnLd6rTA1Ci27Is8sYWt6j+o7uVDApn7HyHWZtT5LKlmD8PcnNHstIC+SnQNyOR2lUQRtPy4y
s76ENBK096/gY2US6nW2GZ8FEVejQWmyi7yPyskGa9of4l+J1JbM1GfJ6+hkgF0vYtQ+6gOVwt3H
mR7Q1b9lLFCEtexr7h0YKYR45ZMe5cexbmXH4sNMkbnI7MTRBLm3QCxVd+/GxH5+CdDImtIw9yP1
JfeJsqfN6Q1BFsD8DAd9aZpQ5lQJQtzg19H2BmxEhlclbcpiEZjDcZYONZbPnyF71IiLMltSQrJ6
EpCBPKMOp7Lp/rxsee6u2zx1grkuJj3fWAiGVHK9knLFSqRxOSxkmYvhOpQCcUAG4CYbxV/GeyOR
blHEx9JfwkzBeppuR3m3Hn9g+x3o5uRfBis+e8pSNJcD8tQ0RmuqRQ6Gs3dqxCzPjKyztdt9d8s1
8X5V/8s2gJ0AYDit6WsWoCY+jp8mQiQPyxQtInWx3WLXmZ+YGOzA6rHGH7X/e57X4XMv65s3aAw7
IgyGIOSnDfbL7z5kZFDk1xIXVwdQwAP3MmZWayxonLzlykXLFSm92CaOK0biSVwXGHfXGwFQPNHN
s9zL7oS+jUp9pNIqk7ab7x32sTPu0BVKeQU7JRjQdWPtXp+27gu91m+JOaWtQ0ioddlc41Qdochg
HWxAEKXzMdqcPmUiKYYS3gBcJ/zjuW4RHgdnOQrsjsgRfcMDOFYd/3rfKX/zIHrydVQJRbSfLVil
hifBg3kirPpws9STBrOKoXBMh5hR+FRLOaRRnmbQRU1DyllcnRxTuJ5ByQQogW5qlqoSelQlgjjq
vVv695AnPVMiMQHhjiL9FgjmnOKUeetRRift7MQNMrKx7kIYn6cfGmU/vfcyWfxYqqzwIMLE6auD
hY6kHfWeaWNvNzDGrZgt0wlpWYCnPZMzE9dSgBuqQh6IJH9OjTbfclYer0JKgf9KQj3nHKds0MLq
6oi7aTdUP3VVTzuIwvu/0b5fcnLxQpICeNQxEAbAo+zzxZsCS6zbPB01Vr6NJL/PZw27eSIBrtjJ
txDFsns6ZJnnmcjR+eW/9ldW2eCw3cCyomHuC3G3pXaZb3C+pc26UajPMzl/ztvuUWtyAAn8jNep
5DeZ2A1G4QMAdpvbrNPs/TQmjQoANSpZaEMTidCZKA7bHPhFaSG1dHIYuIaacAqQ54uX8fJ8QivN
pTEqDpvzJzUge6AVbgE/z+K4K8hjI70SizgXMoaEv97BcBc639JjJVgTmsosA5LJibL0Dmtum63L
6njaSb7KA+E+36uqv9N9g+yZzykAKGAWsjYdoTR5K2+CZjrJ99Ysktts7KO3IrDCyLoNEw0rP8QW
bi4QpXdKhcO8KH3UhBkl9WbWemmicYzT7dAlroMdf+AKIgoOPv5LIJo48NQVohsIgZv76ovifspx
yiH2Dq0dWDnZQOo3i4pinUN3tGnubs7FJsBHIoVJruOLIXV3E70sD4A6YagbkWr03ujZ9+uJR9/Q
8U4Nviz30VXJTKxQs0ZFWxwjnYsOLqGDAEGQ36u/oF7ZWjFUxNuXQIsiyPcjmtHxKD628YFww15Z
zcPHsz8oPzlR9CYKRv5fsg7AU1uThv2ACCCZseQJ/IStR6yWe7u2clmgha+lV+PVeZTQdB/01Xrr
IVHjNkbbVBziDztDI5gMxyytcgUeWebx1PaLwMHLhSeepUomCGEllH/yyiP9gN1Gc2twdFNpv4jl
25sd5nqfGFCkQ/+ikdaeY+SeJyy6gMi+Y+aH4HXh7zXsBQ77PpgqrhDxMIjocPknfs+n6N6O6ReH
gdztcCOF8TS54q6i0rG0txOwRz1pbonHzS0lE6rK0uU96UwvDNPkJHeRwdY52FDAe9VCddSJ5jd/
1jBFzb+FmfFJ8oN/8Kza92h/nWiZb9vci5fwmt3NRj1WpVGSmamHCDuPUR6T6v9KIVWdvxEMyw1l
hOhkulnmpbsabGAIfn0hK/KYJ+bnaG+bCF1/WyFL9zH+f9bD16RAJXPTF9jajQE8HV/nGkp4Yclr
MVocK/yNJcNMwnPJujLEf9rxcZcCBk+zbivdgIsFcug6Vtf5eBFMA72a10PL82Jlemu/k2kAadvE
EMUFxImeyKhiX8LRYw60tN5TFK48Mp4LYezcZy1WoQSbkmpx308P6kwaOB/HSfgtygblUaK1JRuT
iXZNQluYJ6hoY2ZzIZRald8HHspjmwxH0qNViHwqQnlZ3aKKa+DqPefInaQiDvrHyJJP5fpQ/iwY
6bx9r1RbeE8sybuvjXZf54cEd5Lye+dMUItshkg49CavccZX1gU7jtFZAWjC1JpFosZSF/zHdqdc
nV3YYldRs1EMH0nSzqhDp4+NTCQL6qi7dCBI6woutxBIJ6YRk7B2Lb/B5R0vYIxKuSM/FdABIEtl
MFOl7lvvh1mBQgFpjnavdxkZ0jw87zkZdGyZASYpIA6DqbxsRr0P0fWbcZ1LYJtekT8II+0cNT0b
uLl3Q1X1uthh+q2m+kAMyugaVPRy6aCAzyqFPor6OIi+pxnwGYguYupxai/TLsoJ8MKCXCy3D9m/
0R4gHkfcAUleSLHWSugIOJqDZup/tZ/X/wt7YWeH0b1AQN0n8/hLYAsPBEHFcdW/ZQqGlPW+IZiV
zH07W6GCboq1isVm+OncWS8N48Rgc4gB7aDS9YhqzA3XZDIGFvCDmXARYMifDSTzAcFeJzvQLm4r
ywHLr9kiu9qFC/QEmCIZH4ILaJwmUbc3WDppv8BNpHf+1UvuGXD6/9aiMae2pboax/MSdOz9Gd4K
LVMzszGfblw7iyX8M9D0LQZdNevLwM6C9bHFPOJ2teseHk5K2kh42em49aGiG35mU0AsUwzH25YU
NeFlsqHH2SRUBjC97e3FkohkOPPd+K0C49PnesRooltFeAUscBRsfAcZxEEH7jt7EGQn7tRKR/cv
epuo6g6pYDtrPUYmCHikP5GGPxE+M6XeIfjWZemY1O5h2hv1rC/JfiHGR6m4TSVc4fy/LWHjR1BF
uYL+BykDsvdVXF6E7dtbDxBGXIQ1Gb/F0keCIHI6cJN9DB7V07uELv5cejUiYV4V4qycIcLGKlpj
EyNN8OXgxaGX6kC3koWu64PjJ4VwL1vVOT8maBej6In5a4K/oz/TF3Qihm3KFX0rn8i5LDXONOyA
J2GyP0lgYIqy7THU1rZFGuHzHAjWM5W7n4PLLyH5/Pr49Vk4sBIEScD372VJh7F8jcllsjUbZz6R
sG1p8tU9XC6rBRukX1VEseL0PS7sf4Bw0QKiGfenkFep+WtyRGk7yMs6MP75CDu9MdJDrhRQlQUO
lnTBij4Zet4YcgkrVoXdTvFwOVLcim6H9pw5MADbpwutQyGemDTj0LCzA71fERld1l2eZ1XlD0qB
rEo7l7x9xJpb4Zzdww4sv5poBS6eHk+WlSE4ixshVpgGeqGp5chc1dBHtmROAi3E2Cfsx3ObK/OE
pZ+7gEJTfyHlgvkOSLwJiyMucV29i6YDltKbA6BvAKk8M0S8j9XVDUrkFAegfuzeMKgtmOUU42wF
5Hw9on/webt0uVjB0TVch2k6YSV70NIR1XCOMtfnEyzXgUpAb+vDwwhQ+djo6fSahKHJOiIT7hPo
QShdRm9YsYpaViXxsSfiQZvQNqG1kJIQh0P3rQTCmWOlLm83g3+XCNiEvmeLy4NkgIwUDPE/an2m
Vj6xpK0zLll323sMsbNg+rTv9yHddVRCum5HvKgGMi7IIh2WgAjhIfJeOmUavZpDxg2SIkP+vHie
B4KPAM66yZNqgE3dQPc4MOal/Y/GZniBmedyfKkodAVOXjEMYWm/iSocx9mvyk0Va4ZFtbw+ESQy
TnEoBudcL7HSFSvEtwxiUlg+Cjuffa1jHEijLiNhvDlOT6YAU8dbap1rI46JtuUD2DocPNmixWs+
t2cF9BTLldTfo0Sv6Rut6IS7zfvB/PmRB2hFDHmgNHyx5Bz6H/i0x77x+IyE0JdJ0Z2CyDmwqOCs
y3DDc4TnF6up8H81THyJoYIpdk8rvtc1rGN9qGxGLmQWJzam+b3lvuUqzHoulTSK/scXKdnKroYb
YpzhBtcZvwRxB+ZceAu5DtAR4QZIR2QQ97X8svkiOj7NgDj7DLdgmVf40ixvrosLvQTIOijbfDN9
ZHgL17fGamD6gnh5FTSsJGThnskPh2p9e5cQ1ai+RG1G+PACEfnqXh7jAqMr5RwW5nmf5fXYJCN/
dzIVYe9e2lFakDfsXkCAMgVyzmvf2DxYfsFOJDR2DPbMhn8iPX9PmZ9MxtKsuhc+9rjjH2ILrT8p
OJnrWEbjNkeIM2cbOXJWcxk73dxuW2TKcr/dPg2gBQvgmBxrc2sMoSk8VdNBCIbaJ65SHIDAAoXM
Qg+t8hBBVG6OlezoNsoH/XTmRAyt+Ktfi7qfJ2Tx9saqD96qw8gqbtPU5Tw5Gw8vyk9Rjml4GP50
1AIoq9LAqEcfkrSKQpk4sjb4KMKLrwRkg/tXTp/6oNz1wRaoVnqgkDH1lfwDDkQNHARjh56edn9J
SNdfJtOpgzO2ZOvCCeck0wK/8iC4SZ1cYJejP/tR/dwVawOeTX8NBnfhhmW0v539AkgcFeJVHeV+
4OcpEIIupLnCm9IykK6yMy6wEUeJF+FVOjK/eOKldD5PF+cLZYQCEYjctadyBFfIh11bZWHwEB8L
BBGVTUQYRl7jqu2t5j9HApPCopw7NY2u4s6R4iCVY2UEVk60cm7BnUuVq/fpweLBnMH898UdN2Jy
IIP2dDWvHr18WTWViaoqiI65Vo7W0MhleSmGvBYeQik90JgX/A3fGewXd9qODO6dtgNBWjP3vx2S
vB590Hao3RLfTmXszYIIa8829SJf+T8kUVDNp3m0dX+/4sEeENnFM7ARIS3aDTIpQkRu8x/wunqJ
6EH+GQN/AAnHAEzvO92EP8JLFXOtgTYjv2u22nQQyxQRU2KDDuYtBbjyQR4ByDkHc8g8DXKBj+57
bFCxgwEp0PBfgqLB1LdVyT82pIs5XB0Y7BCJY5C2DIlqlgee9dP+k0uuuJxNHz9hMv5Aq5+l+aDt
8/6iMh3jWXxxtXXtrt9htztwEfITFeJolWLEHrs8wcQQFvwhrD9FpN/Yb5HSPwmSFQUUCAxjXHdn
IFX9N/yXawd9Eb/Xp8HO7PyqRuUkw5aN5zB/UWuSi9r+UeD8LgrVD1mgPJWpD74zQRnQcPeoGysF
VEdjxQS3rlrNjrvegE4MvLxYDGirN9XV5JrKrtKnmgelNGxPDDXO3by3u4SpDnYufqUImKc3YSum
Gt4OJ89R8pvDQYcO8v/sFnFOoclkw+5COZBBLTznGavFxs89UxG+YZiByHk7S4YqhaTGhbq3HJfp
+NeQyJLLlnpIGgV8QkjKJ08sWB1RT1Vz9+6jSU+2i47+hlkbIqydFP3Sd/5gLWWHfQ7k+P5CPw8q
F+rSyh5iETeiuio4yqvMcUMdBOTDU2lRYPCqzoLcWkqNJ6TKh08dNLNwvml6T8mzNkNfF0nY8hIU
NrV0gA4aDe/aULBzH19xTE8aY7ccvBpjbGnUoRSzwZnso5QVKAyZrdpEJd3Yi46VmrKO9kV0dp7/
kpCiqfBLqZukHur/+5hqWcjNEvUBaB/6uN4nBvVSjy6IjIdZ5yK8LhzBUMhcILFTqEVBFkD3VIHS
socLMU9REU6bbh/8j7T71XcVULIqzeYKMiI9jxRfYIzj1LRQPLWZgPrx2mOCgLsjyKyPv1slZScn
HYBWGR/GX35i3lb9xYuG6HQ6iCTlqW1jMZg6NT4GPaWCuw5bt9h5EDh8Dz9kV2qfxHy/0kvnujK0
sdn/shMmGG8fJ7Skva1i2mTzwrUJB9KGk7Q3jyzCIkMNQefzpU4125oPRlvyfPDFtMBoYNdEa4Lw
dEPSLy08LuRcHJGGwtzoufLxHDr33xtMDJir2w4QA/Epg9Np13GRA/29rmYeoYvFNoFALj+52ky7
czbDQ98q31LWG3wCHUNIluQQNLqMIjM8OT8BbObRhfobrai7N4jUC0CSyNbXysc+0hhTW/iAyseE
MvhHWjw+kMM/CiK37ntfHZ0UCx3fDl/Wp0W6pUvu+B13WZY42xTbvIAORIZ9+u17jLTphdy4IsJ4
6ErN4Ut6PFcTuBVmJ/MPBmQHzoBdEBT+//nR7cL0/6XdPPLPqII5s/5urZrixfgNXQOx+8hysKf7
tx7x4I4JvpWC64HJ6ZLmnoy+CNMmMtBKbX9D5Vddht/K0duhCp96pMF06+2VOnY/mp9LLuDzyn+q
UaHGUoXXLUhrXTHP/TEPJtpFgI3mHYbIipUuCoDkC6rZ/e3QrZpKpQp2nIzP7wp/vAh8Zpp6oQFI
1kQcAPVWlIfOWDo6I5xXABjYBA0XSf4YZQM+sfMI3o/nRNlywSVW9J2ytz/5tpdgjcn5wN5CcRQl
acIQ2L4LCskhb14RsfNw43dpyAHgq3yTNPjiX/i2P+lu5gLt1A4CrD5p98xiNpmw5k4o7oK2IdjK
Qcp77w8d0hAenkXiWnHK7ubfPLbDYxo3jqHcE/68YK5AW8D2pI9viky4KP3tK1DGyi+nge98+KWd
AaZEBjlMqnLmXaaScnbXY7XL9YsnhG0+VoMSXW/vfJVHmilMZ17g5n1wpWNTzSYjE+WaQIvMeVWL
QAzPc8PpPR05RpMSLbieLIW/RUBbWC6s0/XJg3qxvW9b6lZTpAevbuVqyzR7z9XEMRdPd5/l0T+G
SIw3nhQg38d3zZhrUbvqEdiz3QRNA72uFZQ637s/aFihK3Sd1SUpWS7O91cPzNGaNxT86ddnx6XV
r98HwANL0ed50PItnyAfWD7SglogLOlWAuaDdunJSfshUfc5Kysv1DfEazN+uewsox702mumwIQ7
7k3xlaeeIm4gHOPwvkayNkGmw4h5Dn0Z8xw/hEoPUsPuxapUjW4wD3AAIsofP0aLMSeYGglz53k1
BUaFntn7oH6TbhETqjSprzo+LzuPS78jizeY4mOrq5DjJBqDXoLhNjdAKNI3q2SghbpL3I0QDCV5
18/GgYxa0ElzBMpWVwd4Q7Wgc68u0LU/aPBP+zf1auq1t94CCZ3QW7aiXN/GdkAft27QXDW1Eoca
WK4LyRBpGaNW3IO7WB48WAXIrQN8YkapyASQy+cgg++/b33chM8l6FZ09s9mMuGPJ0hq54TW/6lD
Mc5XW29dIb3vMD5MV44Xq0lNng1mKGvDHSSA/F3JgYCjHy7iw1XF0iuXW3Hl6roeMt4WI90bY1IQ
r7MnZR/EInRTlFLNfM53CAw30VDyJwPfeSnW/1IULbmg7N8yAWGouftwDoa/DHXFdfX3O7BJ7R2e
QjiYHb1Y39o9hJq3eQawRTbS2mMBXsUN5NsxCU8SDGYoWkUCarlZdJ/QxYrmoZeXtqDfIwhHRCU6
TgqLhgWGt2VuyJvEkoMQgvLGgZ5eJVMoV2/7kvUluG42vkMuU4uXe8Ow+71pyLI/kZgv6wnErTIT
dGsehib1RT/IIcXTWM+tRDuP+24WntizyJKpcX448SiE7NSgViCNMX+HxVj81fWWhE/ofj8HcQho
ftjqRtGjMwKPDYjuX9cX1z+B+KAYM49m+L63NTXbggaCykkcwDjjlt4baXY8PHRUxZTZJZ0SnA1T
KXyvO81Gv94tNvxdfM9BbYXC3gZUtYSI/GFhjM1sqQ21RtF3prOgazkFpgGs/9bKuBNO1MCxJQ9E
JHv1UXzRtIGW84GnB6sDE9YgLHyleMSftUtNqBKI59aW45bVsyAJiJa+KnnhD+xb0sJQ3qCMHN0W
Q1wlVb2fmmFyrE3RFkwTl3eO272wtA9HdTSNpcoj9KYMak5rzK6fMdR7f/Wvktpqq8r7jBjwS9Sr
O/4YEv4LoSzNMUrRiRdsP1N+EhevQ+WAMpNbbGPscj/0mdOVvEY26Ej6PYQNlwFowESZZKEhnPhx
NwIjIoDDXnupHsC6wA92P4P1eVo3S6vPPZQynapifgsYEk6nL4x0BBApVVnhHpW7t+1z4YRkSJy8
tvmq+NfPOmpIsRsX8qK/jCQ2GdJmoa3ao/cesjDQIFsY//L/wjv34+Zh8qY8vKKirCUyrK7gAACx
pywvTxJUWN+VVGzL9oCPmDqHdjNNtDzD7J6BZ1wG+PvSpubHHk+/ucMw4xCe/fWgO0CamUhtVpjV
s4I3s7soXDNu5eqLu9yuy0XZgvHIkbUSZvy1pzc5adKE0x49LZlx5bMhRBMAVoR/dU8uOA70m+h1
TTfrd27ianCADXPRssD+7FW65TCsMZ3T6dtduFBAUr3UWxOq2TvVDyDQkNsWZmEGiKCBFZmFUio9
SZiGXCgCvMgAn8mtLOamswPITPTGMQJ0H5LaqYqjm8G5C01uE/UFVM36nVIKS5sQ5lQL4b11jmlT
l2E4tId79Dq7dQFNVNky5FsmhTuq2WEHWMAK/I40gZRJKaLkTfHWhwTRTYa6DvLCv97nNQOc8MIc
eqTZWvDaObZ1QhF3e4XvrJ0oAsP4ZvDIjRsUB/qSSF9vfEG3CHfHtd/Sr2sVXKiaN+u9Upi2G1oY
rhPwWP1hS54SQV1gJKrEz3/q91OQLOp26PoDMWhOX3mSgluwhKKxDas00MNx/uGW1p0+jDpmm/qT
VbN43VXDeFRvvk2YcVmWSreiXhWGpVle+XUof2DAJeMOTFWEH0U1A8ZvIdPK58MGQQF0Oat++bFr
eAZJl94zMFQhhpwgPJJxSA14dBvd6zVJ5EXxA+rymIlemyry5pELKxdrtSgke17U3bh2YPCvkkH3
DQ7/x5HqcEhlwUtIHBSbS3IarNLBAnd4X6uOUxOi8Vr8okh/o1dKq/9d0fc1BI1kFzwFCxow84nU
lb3fWXB+dpuW7EsaoUexWpPfdzTWryHvDAj57HEqd7u7ufBN3lX/84wEC9J83TRLWvsXsqi0GLGN
PRDFoQfam9PNziygytdNVNk4+jBI3tC5SyH70rvd8ZpJmtrauDFOVkU2yfqKozGgaZrULjr+FEwk
y/mGb6Uxf4IhBLvef0nYXNd0GMW0XyQbaLd/yL3pJJbijsmKs/XI+Qa49lBw+a7J0JaDjyvbd9b8
FMKVOyhTSkk87/O7UOUhhTubeReIVl95fx8LcSqSTXnvL+vTp6G+gJh7AbiNIuaTOWUVKquxaQaj
CAM9/Yk1l5GysYvjnfCCVQUNtjsWOEsDn4P8FuhXHsh3hSHXg3nsscq7/hASP1mtZqC/crtFGHsM
83uW/xQPRZAP5FnIF9ZR+HmIA/HKa6cODl2J2JeqPo8xab/4yBeO7+OCqiFfZorRoV70GKa4wA2D
SES2TgG7mtfmdU7rXlogTiVLLXoeYDMULqMPZ0qocSsV53c8dr3pDPV6R0/yXXX//6VfRl7vwnZC
LZJ3puEvmjhrdY5dnApq+8vxKDmXYsGozY52i+Pb0N61EpFCf7z8wJETSrHVeAZJpxDS+DwDUul5
47/nZQYk5KzgEdvMaNthYIftsFU/PgY959bQaCRuXrOyUkzp1IPz9VQqUnqKldxYuGDtiL2zktD3
FFGH34vORnQ/067ERSCErUCnHBcYrbFdTqlmP+XNky5B+cvnlQooCukBFZ82UtbUQwKBTVqKZ2YR
YErc2VW69mCiKkrJqxJcUdt0W4JKL6aBJfKv1/vpLMC/wZA6eS0WwYQjcS80sH6USgQx0tdvPGJn
v8DIV3P1Vfpd9gi9JhAa6UHMqq/sUZKRcIbGioCIsdvUqLLTpTU01n6W/l3jW4ECAr+WEg6zGo2s
kPVAMPSxrzM3ktehwYrrHQvnzy/oI0d2pdb4Ky3d2YV8hPytCvKw0waDfsMcPOOP/M10XtYuL7xZ
MJUhofpsf6TMG5YCp36q5gUBqNr3dfhoPgV4Gak5l+rPkbK3fjIhev/smX6klwBDXtS7+t80PdXl
+nPncXMJ8EiDawhq56So8G+rr0oue0GnIHiDah4zrEgXT/pXfdN1J/QGsJMrQEo5gnVOdtT55pPo
Gue40TO7ONTjUJAoRel0MpMIF03dZNBmb0CqwgR64evOdCiiGSPe19wzFDihN7vz/3DP7vcXd5Dk
mBvJr4rTiC1ok8a72ntwyhySy/hKUQDViWCR7yF6dZ4P0+fLwWxA06IBG/X9Lc44Odt0/7DhR+Sh
8egntDKMiIrCHpQ3gaMVeYWDVB3m7uH27+fyTt4wKT1ixn7UtrfJnLETrLaIZEwHE0MuR7j/Ky41
Q7fA2a4p1xGLeoeKKUrMadDqJQPoNREESillEJjGSASQbyIyE8kTo70EyyDpMxUl9UG+zJM0T/Za
N59X3DhB+BVnFWEkw0xylVQyk+r71qpNqNSspko284p/4dXhRqKVSsO6UvTnta8ouZPcszhOOu5T
tZUtmpULjTS/Ls5thZa3vUbQ6M4A8L3kvxMXABw/GqQO13KGQwbNc40hBQ0u7ANxDaGzcgpebCeT
UwuE4sq9AeZyjFfL4ToAvWdXwFFiItkqfAURFnhUJihNHiYyVMxN1buFEJGOuNRvN8Ezm86nVt2k
9ItchDgGYjmviMhzoX22aJwYhjPTatOcowGXRrTXmCLYVssiR0pzXucQstNWS65bMX+PuOGJ/oyg
WAMhvReF8vwKlBJZoD09cY6ff2Ow7Xs6frwJYEOLhNVpMeUPKJWbwpRzNVId4NT/dPAU0p+Y6F8l
KoVhppyBJmgWuFodRkPgrxKkGIcvzmXFNfrtOUlvT1vOaZaEFV7kRSOkVrTbS7B07ZWO2Y4H+WEa
nrInSas1tDsXYzt1pb4Um5bG8DmM9oyLeD5vdv/PzK9ycPJm64sQr69VIYckr2P4fmN++n/ntQUX
uZp97a974EMIy4x5VKBpCv7VogJlQ5EGcP8cE5SA4QArv3ZcO4q5V0It/q3gqAeyT03tWo6s11dN
HSZ1MbyAgrlTG5AEzg8qVgSucynh4bz4V/XejhMn2jIUbDpTz3JuysS9duvy+0TrE8B5/zH5Y31l
CDt+cDlATLgn4zR5CYsCWC6LyacslHFa9Yk8bWUYbfzwxk4qyOkRE153cw8Q/8PBN1m4OC08U7GZ
brknYo+Y1yWzgh3tw4ohJYtQh/u2Zl4GW6aHGEoxRZdh28gDis5xjG7kVPyT/YMQ7p/jbCK7jh4u
UTSy4x3y96GktFc25ampyqyy2xMpCuw39AkyxrSpjvdveWDaS5aF+MNUj76T81OcSTrRM0WouwiO
qf8FC1T+SBOBNTQ33w5LPf6rgrhmv6VVYxy9q7/nxqSpfnpOoOSqMJzViMoeBqDamlQw9WVv+1Dg
oiZ8Ek7d8l5UleAA6LteT4QonPoO8h1r/o8uv7OwoYycqqSeFyZNdozCim8SKtpeoP3973MFDDGT
FgOOD6bTbmr/0c4O1RSoJdUv4ccr3MBCJcyliRWWvbrS27TdHwlbpBsFD4WoGG+N1c2DY7iccshX
dN+aBpccs/yjbFb+1aFAh4czArik1WyFIMRMwMt0KHjSovAp+Q7l6DkafM6sBie/89cQgI6ibEpk
ZMlLP8DS4Z/nWbvzAn4KHIv+xS+o4s4At9opSoPeq8f3j22aoInFGJDy7EkT5VLPsrOpVjGisyQp
JhR1LFpaRuLWJH3e5SdD+6EsYHzz3XRMUkIIkPcq5NGsMdDKt7Z442hVrM+ULoewxFcrjTeH4+Ov
WuBlpdoStFbpIsGmvtsS2mKYcXtcRSjsmbt+5chrBSRRYxqjj2Rjqb7g7onx4E/jbaOIwtVJsMtC
ZWcNdgYA8Kt2D8pSopvDEfNlWnKSqCdrXRpC6jr9YR59WGTFJTkitTnJREekFRAN/uhKFUNDpPY7
Y88gbdYcOtNcISJVdVDFv2LBuU3+US/ITjRwRzfXYN1hqTSyQrCiDdA9t9qv12ZxyuWTFpEAi9Ol
s+CC4/cFeW7N7UKyfUK8nc4lRgO96dfb4TvJgVXGwnN2d9igDj4gPf5CgUE2geghay4dvNycS2ix
Aom59XIBJXF7MNwJTrmyoesFkYkWHKUILDkG7Tiy+YK95ZsXDBNG9/fLMI7Jx79MWjAlFeDe5MZD
uOyBx7ml51RIGpzzl4B+UKwxvbr/mNZ1JNZo+XSZgj8zxk7b4apfY9tt46rmMleeTJAESuphGdVo
NOCOBx2E1C+hSl2Tyz+cDJOTFyAw6PxyOvCl9U+sPR1oXAzYjw3M3zNYiYgl3vnr+c0nECo5FGcO
kYHxawPK1lVKcUS49BHNKy+5QCW2Ko+sVER6WmeX85NxILvW+l5grXVDIGYqiEiBo4w4saoCBuAm
rbhpWcqPmSLWCAF7Yi8HaqnNZjTy2tS2U2O4j2l5s8FhLNCpDybABJYUrozxzGDXdKJPFv2z7V0d
w3eQjdkI8KmqtiOmmYhLymHmcVqG9BUzrDalqgqNfOp0fXNtTZEOoC/CP0VETOVXmIq7KwBo2vdr
JEuuzhFUvfGSHMQvUUmAKQtre+XE/E55tKQKpjuM8BXTkFKW38VAHuIveWXKxmDRWICJOLZmYr7C
Tb61TRsFfNa28zh79r0TMuLnxkuCbZ3xLZvKRqW2Q4/jGJLu4hD/mQRUCSjwm85L+ZnlNLxncVC5
68bnmvb5JIeOX66/VdmaW1HXSHAG4mU7OpsyICNSlubgrwSYiP3M5R+IcBenS1IZIxBM7RLST9JY
e10eWr9FjWYqcgp1PNhjc5jcfRZwoiHKlC1NdOuJ2fIKGqhCuMPQdmRacl/s8ZyEu1wM/7QZ277t
MSFT+0xYUTfyPzd6nlHTqH/JqYGhVtJ3BkCZQpLR8ZSXfLJIo4ByEhGJOw6B+pgJjv2yVAsXQola
ViVVIjokHzm9fK5U7jnYL0bsS1Q3DMSjcDUTSmsLgVpzmX/AqRKX6SnHhNIcmLL7WXa72KVXXuVc
/qYR//O0mqBTiIXVR2i6GyyhmNEuVIUMPoANF09WjE7azBHJcREktzP7RVBg4rLpuCr429gMk/lH
z9jxlOLnrGrtmE1ay76gvE6C5xVotSQSE1rKZ0reO1kkgRmbe7XRndOTCAUJyaIGLJ1dRjStBiyW
TsIueM0+/7xxei8EVqu19xzjPKed2wLZ/m7G3+IdiJlhsdr7K/JPuROCoEUHyHbd3CWb54voHUu3
Mk7QQYpjdS0xU+p0SgevCG8FGoORkG2jEGwiSUuzbK7s/r57K9lGmPjsWrVRRK/3DfsJEKfJ+C6Y
7YnF2KcPgR8XYvCN6jHtvc6qpFgCZEMudhJwRSuhHrPlOKiMJCsY+TCDI+o8LNXcO6Mbsu07nr2w
pb6VktMD4LxlVTjTgAEuPYNkZFhDvcNLxRb8WO3+I3F3WTjC1glekeTwckYWnMY94ny1vkXE8ts4
MugwLDzEAx1M5kXjK01qgYUy4XbJeG+XYO/YCJFiQOJF4RUPr3dSpGJhQjWhTlOsj9pYQMfvNnBS
OHyOTG5JFk7/z9WXcbW62HJgCn7vahz6mQmZnlYJBcs9ZbR9qJTUGNJunbHbkwCkGzYDz0de0EqM
JkMRJqw+5+NR1f1UCAVaJuYOlO+E1e1e88N3REz5YBS+kW/tvJWL/58VyM7chve76FtPULdrXLKt
ztznmsfLgYodWtdA85Pe4OSuMwBEBRlySjs+ihQlfQbHGVUagbUYxO2GS54yaK06TSvGyKaK+B0p
0u3+rbcmiuRJ8svLcvddamwsFbSNtY/WEJogbyJSLS9oxqM9f/FvDTdZWaX0tW9Aj6Zr7GdzX4D2
AjbTOzCxCpHxhhpv/MIzLwyi9C/gUxn4QyXZJagh1o67yxMvkie09Blb7YsrJVHSBSE3v5hfJFvV
jtMUQr2FJmSHXoYlxLG4162duki7CSAWOAwhdkpf+28kD7yP5xS9mOhV5BW/nquPTeaaUOVtGWuv
2+oBwLJ5TeU6+vMbefUPw+HsBdICqkd8nQllpxLGzjfCBBXpF2Mbn9cDS3X4rHdyE3SrZ6fPPHaF
rPF6/UtiDRb5oDGTN3nlDpczFz95ZC4nyL9ptm8SWYCV2/I2VB51V4g0KZOrE+ZHZWDpwgNbbSWq
2eKrYtryBGpVX8Qt1COdwzlM5psMHcQlaP055rdAxnPskeNj5rOXnD6tooYwi7dI2eoFDu3TwYaf
KaGL3u7+EzlKRW2Ok3NrvW3wi3R20nWsArVGhKWGkAV+ktvoFbjL32b02qol/8asXy/8Ysn77t8f
f1xOpVQfVQeslJEPiTfzoXoZAGMSqKLUrd9z2UZ4Pg0RDyb2xU+8ecbTxYYXAZSK6AbER0+pbxBX
hPTN5xZJZY+zzi70nh09wqpowTDFgPzfYrp35u0Rn6NsGCgQLehYq9ST5WLqieSQElQbXI5v4ZQF
VOvb7NWG5qIDVl2xBivRr9sq2Wb1VkQIKJrs/APrxnTCqzU5L5zYiswdiGsxbA0AgZvvqkKckYn0
461pOP7xfzfMrWFIByqwYzUym9husSmhavwz75KsIAlesasqzZIPKOuoR8BULO385tPbeXSUtVn6
SyWWLaN4WCSHzG6rmR0e9lHhwVeJuwta8toMcz5nGTuqhjl0MUM98gU/M6YHbaOHgZgGfbsITx+K
4wgaLk5pge7DfVqBMdBPbQQJrmSoes+O1leJlHEiO2URF70DDr4EIpeqv7FCMKM4fQ0k21vpo0ef
PKA+yhk1jdSpCgDnCgfC1NmSqjK0AlPgy7kYdZZ9Qmfr7LwPF6m8rUdPKsfooerpVV7OpI8JsoaY
2Nx3OyIVRnrXtdtfsr17l8HS8ekHuaVb0m+VCdW8QecY44oqnx6Et0nz/RwlrWH5t9SYWMJH0qrD
LTVy4RiXld0OwIkNQ4YjrBocUvHKRAC83+Hlw+rDujzNc2//zr51i5fvGCToYXEDQthtJGGrM91g
M+ZTV8K1y6V0HEB1yQ94NInzBdldoCeOsSV/oDRqgcdQ+qG6ccrKOUNWhU7v+tX7GMtp+pE8n1xq
08l/6mvN07+od0L3zGgUKS63W7+IvZEbKnQj0mdh9pr8xj7GLcWpDgkG29kl3HXpjbhkvGrez0NF
YEd2JGPFZUc5QoI6cChiWFNf1uPX7W5Vk3wpEod4qq1h76feZ5nW4MZJL4Q7Ze4nTGmVh7KYNPP5
EBSHuSwxWkupj8JhUdqh0FyNM9kb9YIazLInxmL01+HfjGLA+WDbmDhS9vduOZLZmBodAWGjFK7s
N6zxLUzc/wG7I+jO8IC/WbvVhVWbWtoJaNYNbNG2ZflpkWVAI13XyThdj5YAzhzNA/okPgHJDJ/O
O00YhRQ8apfMsa5dO1aY3b/l1UwbZfwI1CsRvbQNUY8uC3I+vWQZxv/5/Bq0ALZjhugjGNqJGXOu
7mjNuJ1FOH9OMqZtUyrWAIUOzIAt26RR8cPhc0aczba/w0Ey9FnoEhXoACxk2sZ/UMQmvvTaEzdY
ejGI3lmMhmkVATKX7T4uZBSL/x2QvVRuHbZeD9wJeGW+/zzvEbsSbDXcmlyAwmc4GaIsM1rxy7YG
DKa4fmV0e6DksnS1sanhIGGswrRKaa2Bo342z6MIO8tWq7xSSVUN0uw0kfBkOv7pbo5hOGO8PTbm
ibYidKa5xv/Q0KhVwfoB6zGnyyxIWBc8CZfEwZDfWgNVre4MOEVi3dwfLHIdLVQgR7LGiqS9SAf8
4HhITX1SzzeLndxYyxzpyVecJBccyXV8ndxMP+eqVAptZT/j3irsoZRw4zXuE/NDnunueFSBmsne
bqNlIjvkbjxbEL+9nPlJ3ZDtrn44OypjF2/4UGaP1Q/7F+0hWSRxVjJ04q+41oOQDvqM5RzY7YAp
sQ4Hrojhl0LDQndebB/92NbcgA4+2nOyE3JTi/S74/mvIThfJ8xyzzO+Zztmy0jBo2n1PWmzLLf2
gpYgduNncv48McixAfFU7G6owAir89pg+ntcvLUFfCz1LYY6u1w5LWM39zH1xvWAMaw5atb+SzwX
WDwYOnv1BZefpVmSrOxNym2oTWZfxTeTrZR0/bumN6gTfL65TF9xx4CCkBp+m+Y4+NPke5OXBavo
/wxJ+nyc4J7/VxmKP+I0xgLOxXzl7o3AgawTq4/GGO0NZ2160jqU4+8bUWOZsnaYfUWCp+PJY9Qy
53ARvIHeq5ifhuhXZb3I1sDgAc6wtnhZ/ZwV5ppLRfEH0woAfQZAY99MFJC/9xbm2xK3YjiNLuA9
ycxcBxrwDwbM45mReB+RIz2EPIgSQdO3wXhdAxchMyu05XTE76vPmaz5pY2mVIQDZiaxL1BBnTq0
qZ470wQ1FqnmsRW4oQxlpwgpHj5+833KDmQkZMBAwldJpmeANeXzwULGFiurVvuyY5C6s2Kyo/Le
6JhKEDaOW0yyzu/1QQbIjbmiplnMxOt0TM/iO0GKxFKtFn3B0Q1I2PYYNk/3EG6IwAhduxu9TjRf
7juvA85gIvUq3eHtBwPv5FQps6F3dmalvlH+PlVxGMJ/lLMFlgogFfUo6crJ5p41q5QVwtLWL+ZC
sZZtVhkh/MaIU5uryjwIaKNaMNwLV8f5/xJ3/TzmMcpJ2roDG4GHwIE3gJvWg+w5jemq2eo70hNE
MuLHHbx2yGGqoeMOhPflancYN3K7C1eLAbMcDcBlfaH303uzI1HCZiScAkdTtMTrJ2Mw8s0yN4Vs
582+ZxBG9KLzEJxe1ACjvtETbnfeMfxzMyJ5V7fFESkEfR3FZSj5nU2nxDJICrrW+9lD0dJGZEQq
izleRnf/MDUC04gXTYUPQgfD3R1OD+VqhCFFG/zC/TwAlBXVfjBmm53HlpIsWdCtWxFdvuCnEmfY
gVrDOUnHy7tgo49JIw7FAKzXEVtGaTHN3q0+cOyduxbX1XiWBf4IEQFP0qxEjfV5gHyA0qDtKxqz
chczGN0OYqb9c+F4NA2vtp+DW5ZyyYTIL+zg9o5eKaHTQn70hrJ6GJ03zFb+6zSsHaDY1Ql/mcgw
gQWotZWSb1EAmiw/L3NXO/qA/QdCfJtZGg+1dZr0/CiCWyOwoeC1sejI//aaoI/GlAM3v/382Nsz
CEHj/IoK0fw9jytySOW2E/mmvqqc7kcwnfGzju2nabovmakfDuRk0jjXMspffqmVQHMEwpP/hGS6
QGFG1hrq3mL5AGtUAkaElhMFKsur6Lzme5jlNmwN/3PjrhozNbnecqDfaI6VSdz3WPrYidFV/t8L
GqU8HtcLifsEmb7AqlmHsBFePppikVIhFoYJL083axuRITDiAxt3bHyOWMU/5STXTDHfaEHQW0Cs
1sEUk1OWeK//g0LUeH0bNOXiogA3tGEJp10gD4SP70rkThK1sFjMbCAmQ4H2RJLLqCiOHCoUmaL5
V7hrxv+py++e7EqR/S6KlaZ495zhRgiPP7x14BXmT45dldZA6E3n5Wg+hEFfvgmqMHoZnrrD64G4
7A47YQ+m4+rb90UhRHWBQQ2nVFG99fF41dBE/k4XyQUtcNcJCN+oWON2Wt+dXsovi1ddI6zGcW1y
r3bZnBOJSjx7wAsU599UUJbg3c3l7qnGL4KXB/PqeBnLBIfkMmFpG6MMxKcE39uEXAg9vg6Oe+Lq
PYGb+jJWUbKJ45yJaoNb4Jv8JQTnKseB2F7uETRgVZbh0lDtn87x8Ob49e0sxJHcvUh0umdTrgmN
QcmVGb4N/gXbmi5Qtl/VsnTnmyl816Fo28wgETCPbdXqxcd7TKgc6iJvxpR//FIIvpPovK7XJ1ff
WQY65pjzVTE+S9BO6FItVKRFDfJI+RdOivvd6c6iM5P8PxDOFLqqK0zfi1qfFItTzHPDa99jDjHh
c96jAOaEYLNThjRpdaMFd3R6guCVRq/yp95U364UxwQUrJfwzgKGzkxri+woRkTESWsUjgXccdEM
nw6lmkRhbzU95SoZe+8VrmhGHcKp/9gyFg6wVpmXHKVGnoX+XQSgbONZqDPiG9EMBHaW/fYGNUKv
kdpIvet8Nk8/+g21yLJfX6uTCW2LM8P434Ea8Z0PnwZJOvEb1PhNjtLpAhHfO0oixcj1IcEgctrx
KAG85JbkP9mT6JPKOHcmYRu5ultbEwYtkb8a67x1IuujeNXzR912f0LZvWXASZ2Y+PXqjRmJ0UA6
dnIAw8DCgQtC8Q7A+Tk4D8ELduN2HXi4TSJb45KmiVWMEfxcUTnh5Nv/EwVttT2NukSrUTn6KBmx
QIhjpzFfvefys/JA3DhvjXPx6xw/qeGfuI0d2OfKQw6aQDb8/Qv14aEmfTQCmJqocR8hJB9IqPcW
qRpwuV9vT8yOsr0aYHdaEV59ZeoUZKa4ZHJS/Y0J6cZ0NOn6uAfc5OGRJ2QViDpHCY8mutNct6Yz
0m+Cfee9GCEP10S0USgaj+6huQtqbQghBH3E3bkJ6yGmDqnYEuuNIZ/B7lXJtzc1RfNJ2EfAMHc6
NyNh/PLI8mGYwLIxjGDReLHadXD0sf/rOdTqKjw1LeCmRuDNJZo6upz8WuGU5QKqoaQrUcD06ZTX
u4WXchgv5KNB8bF0ZJpyAId+UWk24vMd0D6+Dzrvh6dCsmqRrBeYHYsAxKiVl1f0CvRKlDbFO32M
42NyYTjEZ45DSdwjDg3LJn4ObC9OMDe9VLUdFSTxkTyKM4GlOJCGFVKdTDJeVhVgLraAKVumUjx1
sLlN84piPlExDXV79v2tnc9j6NNoFWHIin8PwleAugXSlKvmiOZ7tiD7G+QaD4MlqbeSqbGw6Awa
yfPp87YGX1pgHJxRB156NR1KjMrBNcX5Zj1KpSLDH89dTCg38U9YfE7rOlGE2haRFcaWjzjvAmcr
+G+cC+WzvXmWwl3QVG3lX+DA898Ljx4eSQTjaCNLt04qSMvlaZqZqhqT58wyH2GUjbsVtYagH+qT
uWjno8lBapfVFAwgssAAUR0/GMoO1Srfr9zxWWFPgaE6urVA3KcZRmST9ltskBQSbCRJpKQ5QnQw
3TrhWNUrTHTqgc7vZub5B7kaiBAMqHPFNDWbYRoLcOD6u3ZlhLmxjS+VbcShN2YfTTed6M9lLpd8
cW8+unHso4500P3a/JbVTp5PeecHDPT1nERlJO8LICrAIe7XV5lgiq/OVFJkLi5cQJxsyA2+FQkY
udQTW2PrnKm5broR6Nmgl8iMb/klEl2mZVYysUD4v0Jq9j/yjxHdLO9YOj4a9wr9yAKK1HLsEBRO
EmB5kq8EyjUMTPCaLYohGyWyV/WL9iX37X6LR5AvNkKhtR3jrdK2g4z++Jzy4UbeHDe3/GlytI2E
HIv9kSXwPlhDiX3xs0sVd2CHIpgWQziPutqTRSDa3TKRdc7+IeLYZxHRIl9XKXZ9f5gO3grSXrsU
4FjQIT4gGKjZb8ZZlqBBx6q2i7fHsj/+o5tOM2AAx3UMFMf8SvxPGK1TMeu1jIvjmiq7b7hMcKEt
XP991QroEux5qG4CjJhHAICB+tKjXS2JiPuB2STVMjDECW46J+e4RP8JOhcjcTBHEGNA2iUjZMGs
HdqX2Ogd9xWJcBTsMnJIoIUfHQ6K6KtNOiCX3183QyA8kp+2r7j5AB+jGSLvdmpMmqyYyrXGPnm5
y4uhPV0QrM0u6o8EUjhbZt/vORQ3mdgzJOxx8cYHjxULei660H0NiFtJiZ7GLXcnVyc8ooMkPuPT
AuBbjajJLJG0Djd0RYYRK8XaPftYNiGV7o1TbIO8qzioYysXDnQ3+G0Xy9r5weSSxM+3p1Z0LRv8
Af3R6W1NAItigLslaGiklsnQrMn5DgG/wEY0uVNssj7lBwl2g+nwtMKD1+YinGB/kxLwdZENN9rM
MX4boDwRD8ezXo2VvuAyPiK7l0UtjprUZFLcwDTMo6CC1tTwajDm7AMv3T4pIPLvzJEb+DuwUiGD
maFn4FZhNrQGyVtrYC2AfNJHD79QmEH4nokdhlJcY+ybnbr9O7sNy4IX9O1/8fVHL3PrvEJ8EUEw
NHr6hwRkJPBph2OWnxj3Ri5PWkJJ43XJVzPCCn1hX3vkBwksBsHsLcyeprcAMTJawS8bK+nQuhfU
Nde5SSEPBDMP2SGaXF6kNnJjJAf7IuVw8hhBUmRjeS8fo0MApcCpElReXmrVtuc7eku+0sVhu2fq
CEI5ANMGbmT4UXqbmU+qmL3LgvUwKB8f2RkS/NNVcck5t1RUbHVYNOrMQnJ+/9G1hzv46ah2aZAJ
5Q3gDUBcjJYboCcEiFhZ2W4+ndpWZi+q64rRsj2VvcXEzCroJWitRvHpLMBiW9D+OOblnK8ls/cY
QpGIXtCUtrVQ7ipgG80QXLXuwIh2mzWyhYKhsoMq6QXjPB7Gq6RMS+Wtxdz1FHKsSHlNaLQKxpvp
2RBWLBg5j8ccwjJxZxhs9VGCUU8p6Le/w8ZvoF7EqmvW+ZJ/FiJrgnpWWVWvO8Wc/UuDTnBZDPrv
DY6LZLvCokoPTOl09MzGCmlE6eR8uWthwtC/bmN7fHHkiov+EarhOBFfJdvF06vo+Rff6BnDsLYK
ERqC3bP8CVfRtmjlSy8y1VO+BihjEsy6j52c0zYecC/1DoGbQWI0w1BWYz9D/eotIWZy6KyBma3w
3to2DZDtPAFoSsf5FAewDzNmRJUOpOZi3IJommETGXJoKoVIKmj5xI5KP3WmxMZBimA8i0VgR1NJ
kAM45oBdLrYutlXTNS/QFpABuiUbUH2zoeGwiTGTBrlTy0m8xmxiyPGt3rUbvAWsTWziq6qBxNqn
6t3yYDxp0lCnGQClj5zjyjRtLYx7LRiPe6mnkaduDZjJ40mHW4utWJXXf+gk3tXVyo64XpETZdb0
T+qhtpGKxmAjWyWFHyBdmgJ2GVHQ4/q0+QO7gtS7ZlTeTM72RqN2jCgJjXXUn7dLd4gS24KdPX5B
riWtLtUQD1Ll6C2Z5i+py33+Fy4nxh06ZviCRSO2wlbNbgZWpzPg0BUYU6wV6bqV7wjIBNYRpbTb
HVe3Mv4Ne1qzF4CkrmcAwHJAdzGYJodup+ExYKnmjZ4CjV3+VPOUp3L7qsQ9sIc29hz0P/ixiYbF
rxCn+zA5FXaIxgZ/KHOidYP6pcm91OlL75ZdcD6e0U7+zZOuZiL8GprpXSM+CTX2hCKzOLB3TIqF
abODqKvFAhZtruFKb+Qtwzbdze+KNJVD4EXmLSpZQSzta9vJR+aE/u4mkuA8LA7MW9aipA88QKLV
XB07tHYmSIFpR7Jp4rsHmX9LQ/vB6JwTXCCLVA/TkTmaj2cEVmVr+AfgK7uOz9QySyxBmcuH/M01
sp/fBlwabJuhlGsVES979RbNpAL4BJmq+Fn9LEraDHjyf2DL6qlibatoOoPiegkyt1AZh39Y0oFx
TAhTIcUOgOlknhI0PcHGbNnuB0/zFKDocoFxrksZ64jvBS2l2T6sh0PPIDrgA39vNkmPzL0c3484
hXlXzyHMIFwCJYOwwZ5Dgi2lEqV2RpfmluF0IVihp37i+EH45r3+iL+QpE4qDPCnm3OgUeosOc03
WTncoP5Lfr72PZZg7ojDzRkl1CrnJNBPDUaP3TgNpnI7h/bY9dOXyjr/52Bh49gxiGg2MvZ/wr3J
7rhLfypAlw7HJ9faUFp8RzNQn1wuWlrqkKHhCZoV6aKREq3FbN2zaraatJzv4AcKn1xsWIUGrmsK
jNFja2bMivrjewhEfsqJsp2L/A4RcCsVRpCleVNptMnqBfJjT0fKbQyfHjnwZNymkvTsO0hW+t2X
fzIRFd6w+EfgcdludkLMwL2fLB5n6KfYBIRQYEBFNKL3nHbLnCFmrpvNg66CoEc3vPCTt+jUPl3D
Xv/ErUVZROx12/YxCd+RDXWPei2gtstKQSOcpQK5RNjYUh4XgWDB+Jfn9lSodYM3n5UegGHbYlkr
vNf2FyBNCCOVs1rHx/79ofBJBk609eTnaBNpsgKVQqg2f65IJkBjNeOcI1qvaAzjp+rrEfik3D9M
cZtGDGFPRIoU9XbFst61qM8QvPPVrWItDWrM9kJebpKI2hrO8BCVw7cijdEO1uTu/1GDZYrpyoA7
HKCGfcNsZdvvKTs65cSwEWYdN6Hgvk1wv2F9+fZ8tf1F8u+PzBGJZklNd8XWShoYMtSnYnOVchzc
8CXKGqKHmh2XN6h7TUTRD6Yq6LWS0IftVlqRfJca4Dg3+NhKrADBzPFlmYl09IzlQ58tUN1DE4HB
etCMhHNTAFDRIA3SXCMkeI8lDr9EPsYGX5YccAX15a03LRQTCszCU+0AZhE9a5kZuMNcTvCDYyXM
0OCB56Usns0DuFp0oZrVcQrZt1w3IWw0ORWgJbzkFfXRgPjr9r1OAqqxkoyAIrWbUmsxI1CkLWdR
m/CqjEcGF+5hycj92gLajZlEf1gbcIMKqs2Zwsy7dOa7U+JJ9CgYFWJpfPHeyT+997K55Ehfw8Hk
dHVKOfm6qkosF32luUcneWExZcXht7RrmP2j7jOq2stWZ3d/9Hp2M0zWG/nb6ABHsMujwGS4pb/I
VHHCOvioTBFL5MIJoezTRjz4Tf1+VhCo2svRm8mkzSh2QU4M1/21lSgUKhx83GNtTqeXT8nD+V9P
Ly8bl8xXXXorNA3vaAkMFRmWTWCZRQwBNNFL0R+1tT0MHOiO11sACxUOBV+CiL7sjeAjSa2PwUY+
Pv3bUZ+50iheCAXMW39gvwQmvXVforbnfFcIzzm5ZygKEJZSqPHzhEM54+oMjSrR5PdVn4YoGUwN
i6cJlgD0eesQGpTxA4s+bLHnh36VPtK2cQt0h3T1LaNdxPqzkUc2lqLYQz4qqt5F6v0zCxNqspM0
wwRnS2ID7V0iMjuPjv3IKt6cdS7ADgpkrH6GAfQHJmPuCILhHFDUGJYs8O4fea0ApNU7T4fg6lLT
Pi2KwxwGdObeXgXo9n3VxQkpP7K7lPdhE2/hL1l87+rH3teMdEY48tAh5fe5JdNlTveXyrAkNAQP
XWAFNCBokdXM7wDnRFDcwnyFdQhYWdpCfkQF19YyiUhpuajFtsP+Bn6I+UkI8wwwZ1RdxvzmmI1A
hnxCqFgVsa/PfRnEd4zg7wbqwAEorE9WE+WquN67UR17YUFRkZurpt1DUOis4uthyaZmgLIac8Uo
uJ0h/VXD7BoAe9arNALAA5sAUpbvLbpc0giOk0y6jWHugFA01bXL+tMexrbfYVk0E8SqmEu8nkVj
oizVAvh5LnEKqHT4VpLi0NCBa5bMrFLzhKWnsqt4JEE5ZGcJ4/HfeJnmfVwK8nu+I/TkPdM7ZN0y
beqTq3ySBf5IgZskJS3GS0iD5/u6pI+gR94D3tC/7IqmSPqysBNiBtn3e44oE7v72mLlSVohu4g1
P/Nu8C3nLMZXp3HAIIrrvFnuJiWIgVCUFoqAT/l9RTDl3dMKU6lVqu9tNxabuNuKBRRfJHjzfjDa
J6M/V1UB4GWlw5tgZZwAO+2emutzS4uJKNq+wrbZte6OnFdJMwm8eTUs5jIWZyJ7Wcfe5YvO+qIG
yiyl4xUaloCoaAWf6OrCPKdErG1wIeWpY/Ni/NGWyqThNbFgxGdkLfYWTSsITGthPdEXqH0+3FoM
oGRyVsTcHbrmXPUAPct0YZd0DAPSHAUrbA3X2lhxf4N4u09UzUrLUd78maVL6DwPUXIbNiO4/pvp
ImqtZuH+mvXKs02XxB36dj3sjeD2UhjxWh7uu0HoUMGkt1xdk4zds2rTAxXXHChJmhEx5W9YtYc9
kEg5ykE7s2I03h5sDXY2PxXXmvEw+otBkREq51VzcxE8tBUKsIFCGNmhjgsTPcNC8Atn0f63tzrD
MtOOnS4HQFto0QlbJIOEUX5EtAPzTjuTzsl9P/Ac0/+drKW4CrA9pmQ4UAq0Is5DXi8kwSxQGw+5
57w8xxJxgzbIhOZAQ9TwjU2hmb8oTZkBwflb/VrDmpurIM6UZKJXVUdD8pfKw2R/gX8LEMf3vTYJ
k+XjZGR6zYqFk2fpJiu51iuQ38KIlFBi/2eFwA756whg6DyZ4uTV1JL7Gahn72eLqxazbQ8gWhU4
kO3LX9VY8JfxpjY+A5ReBtnso5GpRVjfgqwk0Wulj61vSAitI/iOoSWy8pj0lkWsvMhE+wR//sYE
IpW0FpEpXcJchASWmwEToZUzGl1auW+HrgY8fRnDl4F+j1uRW2mIvFzm+g0J6AaMAF02x6yLMXjB
iX1YNOgu+2tLnpHdIY+pN7TuJiRGVuSjMmtPmsQh/b7tmcHHlUHHiqlzUoxyE4f7BQYcDQ38jWe5
s8tQjJBqn3f58vVgr766T1SviNpoHD9YLkSFp4cu/c9iTsUAyuRe3pqBIh+iZ5icphBJIBRTQdYw
dygYh7JGmhsrmTkv3pbitOrrFZQSOluis/OeMKaZXeQIccgBwqV2BcC7Jv3z1+PyXxGXQpyOpmDO
ORVGifDvWY3Fu+J71tru5LKo0a4l+fnlLMm1+iWqkQAariCiwm4gMJZ+iVq/Dx7sKXTdmVhlEpgl
qVw7ufAkDmAMcOYjWPBijMjSCXAV7AmcsxRgc3iaYPxPh9Xb4fYpOWBWpB0/eE5/MViK6G+vwdJa
mEgTeLogF91mgMR6SqNyaBpVWPU4DQFrha5oEE5A07pj72/TygKEvCkv+T6T5pVeAQKswiD2wEQV
WOAxD4Em0G3JcSfiV3SOuJPxCq9CJJkM/HnSvepLnWGoD5LvkmXVZw/N4PjfXjxfJJY8zsHYRqez
EONOhZFsIuOVOU8GKBT2E5DCnBk634dTTwt0oLgL9KDAyD+i9lXCJYKOluaAc1xQ9onYWZ5622TI
fAnER6JlQUYEcrSianrBOLI/rti/HonG0e6w6yFW6cJGsG1gccSXI0gldst/QwpKDqblyrlaVZTc
kYvaIaE8dxUylA0PczOc1i+gI8IRKYzQRH3CP35F35eIt5d/tiiV2Qc79R8UvP/0GZXDaBy+ovsP
cx/sn2YgIGF1N60fpbJFtCvJPHtb70fAaoxUMAyKFw9HPNsD3VWpkz04bymyxZTxfbGQpMF4oFJ4
Yz5HWctaAtasHo3FAldoKJV2bLVTnVxw8ZRPZyzhE+UvfmHHnB0tnpYXK11b50fxLMMxPjfPD5fX
Tfqnj1tIN8n3KnE/jNYvOlHbyK+hJIgAiBk4Y3olhWnt0ajJYxoGeY/rWaD8jPIPdRdaH61NH5ng
p6MOsQVaofHTS8/wFIm2xrFjppjw4bGQurAwmWWMDNG1sPo7J2VD+TGDTpjfULNOw5YDnhtwFZdL
iC0KA24IhOgOb9YfT5eLd+tHIiNHTbCoSXLBqj35LtvDICic+vdKJK4tOu79cViEg7FZ/rsftSby
/pmO96cLxQprxKrutfoBz9/8SDpHUvTADYijzPqYKgIjY2LKM8zyyDL3eX+bBkiB0zmGGvR45DdS
uyo2+dnz3k7rDfRI+YT+bqQvCI94tnirzFna6x+1GK0SCBDw7ivyJPm3I2fgASa6uEJJlr9RxcKS
Ds+3xUK2vmVxdUJdO0sWROUhVSn+j/Cl+yex2tN7AKRDxDBXlcezNLL6xJPU8r7yncgu2IH1HnWM
VV2dCYG3dqL6gOBBAji0nR8t1tyMzvqCWHctHYBNDYZgAijcK6JY+ckDYlJrM2szJFmMDwhQcz6C
DVUJ/Oqp1MSnNHAXHbe7S8oJyYu1gW1JddAemMOQCayVoWhPxZGaOkgMHH/U5cax2t+xrP1OHIjs
8jh/H3vbDIQ6xJqAEpnnAsqakjjmgM8s0jVWe8lGfgj24A2IQbnj6rRBs6VbPZEN6h6RxZ02f35q
q7lR4m7zoRsxUH10FgeJ7oMSITGjQNtL4Hn8LlCTMB5OvFDWle95cuLVPTwttgwcafbHfHSv1T8f
ySewtQeUla08kfWAKQDcv2Q+2CF1P0a4QEFKqLRZyfvC6t8CDFWkl0KT4do3CmYBO5KDym4yp/2H
bAwmTYICTKFP7PtRCuxT4yWYYm1+7uO6jryoNx0QLnCA06sIUT4bzU2S4fqcGBM0BlhSx56tPb2B
gf4aqGJsXBPqJBL1vAicfnP82E6eZYMnuVjWqy/jaB264ci9kelhK3XTrt9Bl5VLn7LFqNra59La
cCKZrldpUDHv7umnt4LK/yIgSxFkVAfyk4Wooyx40ABzNK21tFOYkMm6/Vts6PygBTDUzgsPadJ8
cqkEYOAhNiO2RsQWwFr+ykS6zaDQV31tw8HO2kaoFh+fJ1iEQN3ms5vhsVeu9CRlPni6dBck9zkJ
XHturox/sh1OLvgSIqLWkb0benaQwj3HH3B2qOqY6xLmZw/xpNUNiDPbyckAnyJY3I0ldRClupRX
5XxcagchgHXqy/8wlJhWelEGZiPDZnKvFmHxxdcrjY3Hs/wa/RetAtsZYqoZFeiY0J66lXs1wuHG
vuqyZYPe2HolXirzgrdIHne1qgBPGFh8IsTX0zH5Wjs3FueKIl2NE1GNsuEYPjjQZtHMjYXziKkQ
mrS3nj6Z3DrOe7GH9ZBR0XJBdN2xNvTGv93GSNmsGAbT4LZc3HW6hE0y5zn72RxQPi0bIK5LuuOG
swpQwOoTZ/8pTrXmdX1VaeTmH5sBPmpkHva+K36xyrEnuXwbECCGZIdyNdbT3x5NgCOFTv8paAr4
/GLp6tu8FRtWUdwByvHokgVJSQQUOtojroj+UXf8WtMnPCMkMH1xeEtFh7vBEmseacRC8p9weRQZ
l+3FsdBewCzDoZ1QH15XP+RqhFjfGFbDTTdRlyAP+J1i181ZLVxkZYxgjE4yMCCnMXeG7o6dmKiJ
Iy1AfGQHf3HfofWppHKHVbxb3+bKTTo4xxmTKoqbWu6l+hXW7xMWK9+d6L5CkhOKrQmySo5addbB
5HbJsx1iIUyLWN15WNDlh4L+zsqxfD/XVzrASNQDfPhklcrM46Kpd+z9spJn5UokxBpKam9kDvKW
dZT4tRSlyxKNoMHssF9uv5I/UjP5uiplrEi4z2wAbfQF9PpvFG/vNvdv32mRrxCm1Ia1XJmDayqk
qUo7vLgfkkbtYg3dgEohXKIhXnQ9B1FhNvNq9V47HnS90GTknKsRCQDDrSHJeET2D6Q1YvaAG9PC
j/66REUVeBfwKMiM8u46JdVpy7aYQAXnlEwVPIg8UsmHDJDD+Y0a3vCKS29wxjd+QAahGqYay8kA
YCfJbsLuYrXxglM4EZ9kR9QtPJXFLlRItuuthyGRVtbaYQOnMqhuSXLIcauR3XBsn1rk1FeoB7TH
4KXRdc9d0fDE/O0p0begfd06+FNrxelgcbaouq5ixdAmnUXwWqtuZ9+IQ/qUDL7wb5dSAzRPx2aV
kFF6avMXdXHJcNDFxoHZUpoHtBScsZ5ydK6QnxXNTlfZ9p1Pevc6njtfCvsAXQ40io26RYhXTSMr
XE4MoBq9zSJzHtMabusEoNW5W346YIPCrgF0at2vmQ1MOBC1vmc4WvxLUPpLuM7ktj4UWdriHJHX
plj08O4I/SRVEesGYys7qkGSGfJuO13dcHnIfMKT+RkrQ9vBI/TWZjTERFVKmYIsHay/oXa60ic3
NaRaT5K5DTPgv/dWhLAkKc06RzPn4+xyqGYaJRYjrAnNrrFkKmKqSRfYEl1dd7F/ToQjpSBi5yF7
6ZPWZWxuA34aF6LMIwbxpe3OojG3T4xJuFTrBewMZnwaskeMviwTPpC4Qp++mdlT8Y2Y1EIkbMAv
QVkk3b5+15yBvH0mKQdoEOUikAc6DNR9sh2eZygHF7b10Hs2hjZ8ApApQZRmWlixe7hJNVQKhlaN
dXIX4yphqPlZrXk91fomIFP7kY+0ZVEDhN9k+Fk81kVeIrTDv/3Jykyesff29ppFYoW8tOL3V58l
GVKcGf0seqKgOebwypvKiWw28DHhqXyWkurhmRqrgfDk2ywjjnwyu0i4YMt+3ALuvzeNwVy1zxJy
J/1oBdu6JT9vdOsWprcRxAb8K60OeoeacLrBD+yEn6ni6uVJSUAQrlloBTh5GWAk6iO0Hw7muRR3
JHsnn3y1crd9nyg0UKRU1qNSinfogmfvdljvLZBsTDEIWRO4lf2jt1mUUe8LFq5fz8Qws0dnJWUm
GKFBvkTkkdiupOFW6+EnX4wYLGlPYQckQ3bC51G9cmTksmtfhR17tg/AJJkWJA6lrHPcOjSpSO9B
DzDNgARTTgTvL4raUvxMrsBHj/df9Pg1JYgCePhz+Nt5fdXa08MEhmavFU7DecyeYPMS6i97Amzr
Nn+P+OI4rRWk9QuCCjjYZOqJ4wKeuvYNm6IAGoicbOIwHH7vMtpLl8TUnpnWQVgu5KXPV27Tm5E8
COfwos0OD6ozP7D04koBjtx0r2Vm7pBSJA0MmQfLw6P1awpUT1SB60z9my4ePi2x4NjiaxRVJFOh
5H5V3rQsZe8QayHEA7Pu+yWI9OXIoISroKya67S8UgKx6ILLD8hSkNuQU9EKoyRFRAEnJebyc9Bm
ZThyptDaXj/QcLxNLPHLSYPsE/n3LP6woFZNkAC7Z3NFVaWHFVtWSdi0BwczAt9UZumXWLV+b0OQ
Vr1bDLV9VfTB6y+pp3nsJ/+Jdq/74hdQf8z2naMIiiskCCbwkObfkG6FPJQ+a0QSiFQrpjovMhY8
C0Nw7wMl9cP8LnNRfZFBpA90s5khpApWKQRFDRFExMaDAyC4N3m3jRJHmbMmxUWr6TbIkq72VTIY
bN6himhsOTe7QtrmJkp2FfXDXwywAKvCEJYI+jUYn75L81kdQ6ZVAKv3oFJswTuv5d5AeykDpvMK
IfSJt60lsghIaJt0qO/UTM/h9nnVnIRExA2pW25JKyHA0EFn5jp8/xjKa5fjdy+ihg7dvPp1U9ZT
38wuXVItJp4huSaHssvH6CKm5kggr5cV7sbSTzWcri4+L7KQxZ8wPtIZ7uML6pePnzgL/EPtSE51
YdFD/2i4/1X3V6edvDaRydz9Zd5Me61ZT4y2ykX1rw9RGQ7mqP538OydUAxprJvI9csEBS3O3h1G
vHdm/RxJmsBX/B85tmXfFytjBQzyztIAU29trKmdZXPP/DmwKClkgKcTftBtI3f3y2EFuqsXJ+si
Asrt+iDlr5Y+c/L3wJU8+CitLUq2eXVdsj6O3zZTuPZiba+Ayq5/SdE+ImQIKVtXCF9+rlrByb8p
UTG8zJuv2bfISspoQptKYS0mEaHS9EeWjOX4tI5eAa9fRnltVUG8+4OOsDcWIcsK1FjiSu6SaMwp
f9xnrZRb3vwik/3GVhtVX5RZSFglDERH2TzWoap6FY9xcJ+7hfqdmGpE6QEP9dsKWCLYgg63PCmU
nY8go5Tfe3I7+cvaKWbK2kd0k/ndUUU4szdhdXRAjbS5Sn4q3sxO9qEZ7we5AfJubG5njmR5TriA
3woa4dubHJxE9Fj+cX7A5s9GXPxlB6W5tmcwgK9svMzSPndbbLz2OjH1hEFKDFgq7SPu67nnrEL3
z8OrKG2whxUKMb6TneHnNjSvrlwggvqjf6OobE7BcUgi3ePSV6trHJxLnhtSr0YZzL79mr7I46jy
SVbJ/G01uZvRy3VIlZ89LSSNLt7utKHq4cIqgqZzOp8ZV5kkaGQka8cBda9m6Sc56npvFx1+pZty
5FfhCPo9pbRbFT7qAq4PNY3GLo0UfKIKRTYyHOUIGPpQCG9ty5uJa7T13gqEv0rTS/y2ma/trtKm
go7Y0UJnFk3zEeQ2FWEFj/CqvcNDP6z+Gy+5iTYO9V6s4t7tE3yMatp76wfYGFbmTF59FgZ33lc3
e96z/NZRsp9q3YZFaK/rb1N8Q1xGC4Sb7emeBCmrvrzrs9PrNFwGMtpIzpB2yLuAXgyMU6IMJy8x
MIVcZRYZsbMPHK0c2siWLB7AjjeCDHUoNKT+evdKCF/TWWLaCDuQ085AZC5MV5EYWgS5P6Qu+bpL
6uA/kVqmuLSXZtsq4M3q3GvEex7+Qo6W8Lqs+OlTe+8NEKOuYCVk8jEVd+SlXsnCrAbbWIKC4/E9
7Zzv5098RXX5sQcREd8WnG6no8lidIY+JnCGKp1vfD8ohdU6DWWNf4kI8qZ7yhxzqy8JacrL9TPY
Jz+NABdgIFjIfOZEkdiHztQ8ypVkoEHEID4Cyq3sXA/4zhu8G1nADqSn8RkPeFkaw+4s2iC3Hg5x
rOZefkFUYyK3wJFCbGN53dmp7gGsHi9Js6XCCp9NiPCDV7UIPhLmbDtqgMevcxuGSB94I4NQjCld
FiPMKWc50x6hTXnIwiQfS9rgeJ6WqyOTor7ppEfpQkbD6oJh0UQ2mOIYKDxhTU57G52wV5ZNou8n
NW3G3bp6Fi58iKFdJgcxG/V3E2oGmfV6X9M33RCM9KD/woZ5HPXKZl/pONVoOy6obV4PWFWpFpeK
f+b+NBZogPSe3vgrcN4JYZmEaBd7A05y27mz+Pf9S9WHoqzqYwT/UB66p4T9WjCg8sUUoVS/Hi78
IPCvROkr6xt5qkYWFuNXi+PWekSoDsBSplAZgePNiz3beJ9bZoYmbnwMx28Kqh8B9RzasPIHDaHc
fRCdZ2XBY/yBecGZRTwJbzcfNuufJgbnjMw4P07qSUJ/ej9QehrvTMpzhNgiPe9YmQ23Rg2zYX8x
VJPX1u5RvvdPEQtrqq0/bcHeZ4ZVMdGYUNbCxPEbVAjKS3yrRRifD9e9CJIfKxxDsk+85xAS5oKx
YVFCeQzyCJz+gvlMqliau9L8NSScx8cQzKtbKqzu629xrXu8nl6M6M21yTplgVPi04VCS3mg6Zuf
OitJjfahx59TS/T1lqH2ReBYq9hfPLjGDKRNWmGLNAOFbIaUtDq202quKrwZwlKGWSixh2hvpLOD
KZRVVKBC+zszwMLX+9fr7pCDa0iGTlaGlGDNO1w+wFqdCBmhrUP0MsznXTKdBBLKx/aktVaNazFa
JZWDPUwtRnktzPRXgIOdTjdh6Vn+tQuIfVaO7Ioi7fOgjfuYtn+6uQ3FMUX+0T8WA11tsC5FKXUh
iDimSgB4/abaXavtTF4wo4V99UdgEHSqE1g9McxuG9mUylg1ebbtnXubZuTuex1NC/kNEJGw7DPM
NtlwpPRpqWcKYKjE1HBtFIAOBmABhL9YVAoa9EQ9Dgf4yD7C1rQnssAWbYF7Qp6qsUu0KemBUWV+
GE4lhUdNUyCCeFYROpY3i91FaLPIfsr6WJhlSwOlLFd1Nf8yFCE+2gGD8zE1QPSAmgba280RDEpB
tQKjBWXmxXN2qsxVdPJ3Ys84gToiewHU/GY/yq/ex/rKXiYqIOODRDSYW/lMEOVV6F+j0lozVIE5
WPQe2qqfFTC4iVeLhl9V2zymVnEi+1tudemo8HE3EjPgiL6Fn6V8+Eg0Vu4kPd127gnNLe0BShfD
QZG+6p6CRbA2YlzKK1n1QLT+Gnix1bfy+a4+rhFs6+hJWCHwye7UjdQZZCvj+n6HgjQe7NVjRE4P
1FPmLCNV+M1JlASoQcjBthI6+lgVmsgoFHbjLGbJTs/BkAZHVrZQ8XlJ5xlB7c7nRnGUwLAnYqYK
bgEAVdxBsKTsNo1wfFRylix32UoLNPgPABLFOa7PlHURRsgSexHULHmdORJugQMT885kjMd4GEuC
rYtCHv3ssNY2fpYCcgubzP7y4iL3vrr0BXCQEryvMf/Zo4ABEPJOnzvxAW05OGo+ZzrJ1/uGq6SE
KIscwmZl2kpgbJkKp8XRMksnHO1sql9LrA2/4Dh0Mq8u2xIB+0vBrE0kOHC2A+77//5rL3dGvv29
tet60caSALWugaahK7M7BaSQP44FZKNyRJWTddGI9g5bNOehbVafNTZwKL+NowLqHr/ze6GgB/C3
jnLroP8waxIZrp886jePyTt0FsherMdYvB+k0YvTEdBLGcAMzjYeFvSFPddZvC89iMBbReImRKjQ
TIoTnpIBMGDZFsUKoPZntyrw0Oo4pZtVzV6Ayi5CywsG+uFC2oucN/e7fX1yBtIF9W/ZDnCWvLBM
+mOExWHXDT2FxZO3PZnlXHQBajyWq00eGx/1ktDJ1F1RWz+ZgNqa+5TuaNLpS415VcQfYUp3rRWJ
6YU+Re/JKGe2dC2kZBTFBh4T2WPzMs6/YZDnVZQxA3K1nPXz7l7x/f5ReX7y/j5JYg6Qogb6Uq7R
SRos6RLCq8ptcUHAwF6M4p7dk/SQDtsufmFEXq+b4bj+LLJ9My8leiPf6TQhH2yIpXZuxnnU8tAH
5Zci6KoF69/m2WO8yvTMpA9Ai5E4BPrGKgruT6FiklHsB/OZbf+lz7CTy7w29M3RsWdyKl2plPJ6
EaYu/zONgaPk+e2UCqw+H3vJjt6UUITYKsNtGcj3EBvY/JPR69RIX4n/VsfTSeT+KTPCekVJM+9i
yuFaUyP7rN6dzgReG0pDTO3IWXoDkHWW8rYSrjlnzgnKrpGAu4RuG0L9Km0pbjB7SplB8EGqfNLP
J9YLR6gySGN3535nqnAe5ZRo0ozh8LOLW1DMx+5naIQWxjXht2PdTFIO//UGbXBsPncVYOg5nPUf
AV4ODIpX8p0knKz7CAgwqpn6Y5krMAWmf3uKopaZM8FuKO/GJsB3Z1XEyJxX+G1uPvS1bRzJ5tT3
4kHEYSXx0V4FK3ERr+2okeomImWBFsPM+Bdoo+j0CfrjFLb5LSjfjXPan41l9yHftltq8MVcaUau
rSHRJurNHehRszKcdC9sK21qy7aQ/qeWZQw0KafBZr/vBKea8FN0F3VurvS1HVQJs01uHHjfioez
0tmTP4oHg3Jvw2DbRNcR/l9Jft8fHhjqLvelQ2oM6K57cK4tfFLw8o480cAuvabmYbNiUpGAvLkY
ClUdriyleCaPjcF4Wr8kseeeWW5sfrk6lkBEgM5cnLUayIBrU8ITnatUzB2oS3kPgiGn85pqZoUl
Ory9cqvP2ndHpfB529qzrRqyeOWN37/gaoelpXae4rDb+HOikQryBSU1uHP9Si75S7HOA/sWiKBZ
Q494ZLBKjMZP4fku4R9MolYvefQ70ZcMgQn5tR8YFRFNnOL/vAjo16illeppzHx5Kv6m0NzGmX4M
F48H2/b3jpNbP5Ep03NXrLCZ9qpldEPXXZgV2iO8C8Dw5iy+vG/a9PNM8orPXQbqNXZHyUMFzu+i
Akf/zuQ/XLCVNgEcrXHRInmeStB9MeW/DrfJb2EHFmmsgy1IpV3+3gPYF0m7yfyKmTlRxJTm/zyH
axmJyY0FA3oVYwvAYIUEddsbCzgwQntAxgksrKxr1KA70HjJkdVPPVrsPOjXN77FQyvZJoPKnUh5
JEV9MR9zmTNSOhBqqfD5WPxmJ1UxdKGvCGnXtj1xyaCbSAPxAhGXsWFt6MNvfDUyZLZvQueM1tcX
d9Eg3Tyh5ugVMlT8TMuvSDFFqblmhSPl5XMKtyF06tPnoiLGV+l2z7kOk32biQrmT4A2huiOb8o1
p2D3KpTlvzUYpbC393EwoBiWy5dVyBbTLUp/0ftboN/XdwZbmulE4QbRdIgjnLBuEcdD+3+Asmpp
sYo4bpR4g2O4vPQpe0UNf8G71PQ08uUgrKG51h7XPVCTnR7HG6CU8yisxjn6siQRRjeDPtbiss3q
qqDV9auWmrkLk6aVteMMgA3b0vwRAWMEZeWA24xND8spAaakb09TUjN0bt1YlN8C9f10ZYMYaLbn
yEEVi53CEhFc0ZPejyGyqRqBbZQVy04Mknyj0ssoNJzhwfQk4fVQSV6AriCNg/YomiggZ1UPpd1h
YdY8Us0zdqFiTKodbQIzDoZuQe4gAk1wsN7FcZw4rfxw4R1bI7uplvNHObcaKykJT086Vw9e9oPX
wgMA6M88d5VhBYR9zEuGVm+edI5mWM0FTFFah+KL3DZVVOcvuxlwnfp1YpQLWmbWHLLPTDdqlcqi
HZeToDcRy68Z/NrVOLc2izTYVWQsugPeHKtPOBzlsfMEyWlUhKDRkcIL4NlrizWATE87KdimDP8t
gZNZ7VBbL1GGT8tcKl43i9QQG0XGFM8ATn1x5HGhvQ2FYJSTqdI6U/I/j7+wkMyz32QQ2qEJZNlP
bGE5hQGqrMVzOIbGPL1IW5j1r6G/xZru9Ij7g6pZDeRU1cS3j0mLiCEfbjMWEJBefak/76bSkVoA
iW9YKjQ1qSdfLaF+TaHSLDWML+VwAzgucBcQi3sCWXjjllSZYN6FgLzI715U4Z37uLFAlLBDAA4s
5WErR30nng4f3QI8y7A724Ufd79MHdJDKlyjP1RYhoweIJu7XlpYBYw6wpd9BFjIQsoH5hywyAZr
vl/bD0fqEq1CmlANg23g4w2lfH5RLwFZCxPPxlbSXLcADLQB7ooi1+PDdIU2znOA/tKmbggsqDse
ytINPAgd/pwsvGWGIB8zhSfueRyuDMqNXD/3h3OyMvUN3jayJTjNxCKTDEpzXAVlNoMy+69fRBlP
IzCk1TgVGUFeSHR47LFAfj/Y41rszSGmtrSCgLXuAlCl2v+FV9fI7xhFnnlcxkHYWw/fcBejMHpx
ZoMUpmrgUB1oPCeu+xRU5H2TJUNJHhpffcItm/tKdeTCHx3d3sVqn9o4pOfQ6O0NGsVFVF6MOcwk
Pmpz7pUqawjcOjvafsHRcd+2vCOK+W/Pp6OjXUp5S76bqOWU9D6pko6wODpn5dtQKSh8AN5YAhuy
1UosNZank/1Vmjair/AP2XyTzF51tf5C7/WSv2KNIjykLDtHM2dSOcPxM5EnmeMnrzhRSWFWUHOW
OqouwNmTz4D2a1bB8SM3G4vC2sIQ8P5hIBaQDs952eu+CIX5RWP6UXgRG0u4n5eezklRpDKC1H6M
vZ3UHxF28AgCvqi0kXhM170KSBsFLeCRswnhlnHynMmXEp5CBzdJy5ZCRdc0hPyABWbbeDoWyzRI
c1KneE07x1WS7g6uhN2jOiFcqy8RIQtNo/Q/NQ4YEKDxGDGL9VZlNhXkw837+pQvsMpFtdD6dgun
nj3C6l7Lln1fq7DX3RP62owl671Lzsbm4ZmsPnNx/NPLZuH3fGtMsJrCOLzgdRNjVqjUY5Mt41uH
M51q0lyGkx2pITipmcCUGZLZAopM1vl8g6yp9QnqFbE7H+EZcjh1kfeflMMfM+OZoSSHNmN0p/oA
MNTVUkh6Ho5DipqeOKar5wb/0VSRg1xwvaB3v+Yoi8F/5l/Y/9qdjltKmW+XY8dkl5pMGC6pW8sz
yNtc9ADMUBEeala7wAw3BI6lgVR5RCvxBhqZVQfqZz2W5glrOEfeL/p4ZcYKtuoutQMyp54HqkDC
jKaVKPXe94J+6pO3249N8/DlD08UJSij5KZamPHSINfYq3Bt+sHTi/p0DH8EY/OLVsW2XK/MHYeW
WgRkhWWGm2fehaPxQZrN24/2Yj56DPtguYOte22o8PDpH6RzWygNtmIlUIPu6T8dXVox2h6+9A4F
LuSl0OKbe2xu0gCuF6j5rbF4oqKb8sPPSOMIxfkrZYjwKtsaObUFF6ymD+WGl/TXDZFQwNFK5dNK
O2WQ0dRE+HPubONrl3Bk7+81COABq5bZVrbp1JStVtTFzodZP3Bs2K598eff9u4PuY9kLn9R6Nyd
ibSTtr39t3vVEQfm8c1i0fo3nvSVEoLLBP9qKFesSInuKM9zr15DBkzUiqzB5D3almQc637sZWpy
XMXfXc5jBcTi9Iwt+stlTHXOzz6p7Gg1+iWZKPG1SF8oUM4ZdsPvZoVhAxhZ3rABUBLsdRGEQV7/
gnWMGdYgrLBW1Njrvl80MrEpKbpdPFCR4hyn2EaMcevNTBBVi8CuKHnGjoYhvddFcqyDEiX1FW3g
Cszv6iTbhVoEXjQuihAL+43m6VpplPUwf7Ss4HwXRGUCzbuL3QjeD8LXN2jkRqj4XD2kOu2n6jdC
9zfG/7x0l43kucIxsJg2EGS12ueKKsIJ84OCEh7W32QtSI/QcnNwmScdOs1BqKp1nxZ+czyY9x/F
TKgRzvFi3yYYjZtn6Oxi+mLcwMrvc/Ea0bakjyXHmjbK3gvE1MAw3+Ou5bauyKl4b2QVrgdGQFZw
IlbVPwwLkdMFtxI/D3l5CLzpVuYTxTByVKF70RxCCfaqM0CuSCV6wdkrHdeG6r1563y1iVwv0u0T
o9cK3L02J1rIRPX6ytdcksWulNn6c/EvisCH1YHtu0xuxOijXqxtDeLBqgX9rnMH2FDyY+afbYYC
d+NxX+AZpbglUneSbk9s/R95ZXLDqrVsP7IGGZO7khQF8bw6+0bMGXkNG9XBLXxOYUBq4J2DVImh
lc1uhL0kVU+7ZnoGnACrqpyHTBa1+Ofy5HComIgTbvJ1rdA/htVBiJDnC4gJspxy8esRHsG+Q9UT
+9+B7Xr/VajpZZmOOwqWKY1Hn/0U1ccI/ncXSJMS6uek0aADJ8w9TirwxPzboNWLK35/jLerDm5W
efEXQbFumUrD39Rsu/o0ZKTQJy01xHx5PfNG2EmiwhimQ64+nxznNRoWDwX08LoMLME+YemsMQBY
y4RQGA7YgTFf71PtPk5aLBSLONIKmbWrYkrMCMTiHG9eHhI/xrNjo+v1ncG11fOPxTw3MyaN2RuF
fpvY2ZQx02s13AN1j2pyskvNPOtBGxtZ+HzalbKof2LbFaAhAT0E9c7taijuEAZ76kTrg7eYtSn6
nBPrsk//q2HSoUf9F2aA31WreaEm38yxOCS8G3ZyhNdp62mtjQpok3RwSckZDPxs4aR/a1QdlkeL
kGI+xJWPLsqjvamgSPfvuypKwGGskx6FF+sW4F7w5bk8qBoe3DWHfaAvac0juQrGJ4KTKdL2AZpx
C4oJbjPM1s09x0u5K72tyJU4Cz7qRL2vxZBm0FvxiIC9Oqer7djrkpIelTrqp3Bt0gS36Si+N5pL
0/d3nJtn+P4zdtxhpXCqyNyaesC0QCuuiIlw9DFzCweASdkw65n/MfdvbENJzEMKpck3wd33GUL7
WxVoSjirBLB3t6itiDarvTdI9pOesDm+afe+uKw6qcX3ZKPIE7i4rxU/cbZ5j4EyWpgyFQW/7Nf+
79RONakBoZMT1maWy0aDfAXxUF/MwszWetBPBZEDOVjjtdu3+GdN2TrSrVLCmLZ5Ca1w98h3w1F3
/kO+aT9B6lvel1pGedTtaEH4yxdXIMlmsBMw53aTJnDJ/0rptbunv6YlVfjSl+vlYOG2mrBqn3tj
K2bJ8bWNc7mUyhS3qwKysxtOAMqaIuL1FScQRTRsyQSZM/VvKFAwTEJsmRhfF9P3X9DR8eTtphu4
Syg5zBeJ9n66xB8HaOAZY3tKsddkHcTZvejPiEb7tHSI5eLVG8qVJO6+nOuD4ktlpsIA2cCtMGSr
q3u29FlT3gG3vyiC7HYlImS0Hz0TBYUHadfbTBrYJrVhQFvh9wmCG6xFTvV/y/YY8B72EfLWlSoM
B4MDsYAOn/BArTHQoq9zI5GOKtS37FGoxZ7LFDyHmhrHiqZj1dEKrUPdaoejOBulSbviYZbQYvjR
SwuE/MHupXKtC4tYlU3UGEhVnls3V8FJJY50eSqYeoDyNIJcIeeki0mmTsVikjOX5N8jL40z9ULj
mcJsOAbfayFIzFGmIbBnrKEIsKjNavCdPCl6C4h+2gtBdjprQYvCX13beP1ua9rwnrkm1AsQqbzC
WkToUqYFXjkoPBqigDGfix817f4VfH2dAOp/WqtkRpgrUwMtfBq1Ur9Lc+wdHQtILpa86f5/UF/f
GB6h1OFkaOZGSZyic84tBhDkIq/EJm++Yy4L8hoWq0exHiilnuosxvhT3jq7tW0tyXdm7clZdW1G
bW9AjmvOhgYkS4/SUu5/hB8sS7B1/px/RN/TXSnbZUiUxufpJj7QF+AAxPPWCsn5EjjohfnQQsOQ
lJwQTfGbNbR1yRcILd+ZmIpFP5T/WH8yK5QT8SRPnV9UAl/R887TsJjxbWAXW/nSqbKy+9rOnYYA
Q/hSMczb0AHEfBwfVTp/GbzkEvwX2yDKcOmR5jhzScrSAIyZbCjiPWCW/AcHnUL3sAX4Yh4xjDLF
LH28Nv9U9AoCuKOzvHr5v3dv49kXEjMtWnVgi/wEsdYsqD3h4gzI7XRfdIoKM+1KmPwJtMT1VSrc
PJSlA1ZkrEQrtoGgv3B+ftkachqgVQXA6gOslj1EPB8481d7hAC2gX8ngSyTfpD44PLUJsJ1bW69
X+9nyVHw7eEOtk2NluQbe8ZoeOBF1INVyFOiS5MW7D50o2KA1vn3UsEa6XMIL6wTABYbcP/G01CF
oSwHn0YHnDRx6O0K4zDujFe77c++bU2h4SrJgYlk1lP16KqkNP33AKTP1DFTqeW5PKG5JTEFLEBa
WY16pzdOYxzVFR1BLcJ8IzDgjEARejf10d6UjXrTAR4dwbBZu31S9O52PhuzrLPWtTEjLCRgVl4w
hQRcxxxyA/32oTuVKUvo7YPJrF1woHr95GzkMtJSkRWFxrTCWHPumePQ0VP61unxcEIDgCTc9g98
gaPpyTUvnY/X/DtnNpy9QEdvBswpcfjaBuk/+DBncs4uAU9UxIB8ZUwmJfiYGgkoAY4hSRMmDkIP
eY/T3XpZ28Y88PDkTe7bOVKNYfGOOUa1uxMu1tpCQXtWvaBn73uug+jSvXJozbHtQ1bku+EZNV/i
GVwH9mrvwUvoPYupf2+zBBowXmOy4VTTcTINz+ePY6fOuZgLP2qGrbfjDW+J5qX8DVipoL9TDFYW
6LhlgE7YhaqbttnZ2s/lgJqupZjWq6wm3EuCtJs2AQQnoLbZrhSjcI/u9pXIdv4FL8r/VP6hcDpk
Rns60HTD7EKNkMsgOZcHjr8lxf5A4+VpSAhSYAzHkIgqKBex4wJNYxrAziKDIj3bZkxp62vVBTcB
TsHS3u5u5pJmcBH3HAV0aOh7yN+q7vDamZY3hYxOBdOzncDkgBEOSP8Vm1scBFp8yluTvEhdeWc7
37GgYyrItj2fA7t5teLI2Nyb1Yskg3j4dNtfAprhahmv4z3FLMBggsjkK7Ozvstv+7S0Qqi5XGjE
xxfHqV+YkFqETz1sVQWW/jessDEls7oK7MDUF9trWe5NtqH1v3/i1lXi8sdZIF9SRj5bOI8vRrJX
5/QKVrrJDVVpdDTfBoZHXPp8j0bdXc2eKIqvS47S6ofAtpM6oVtsZ+6rdAtXZcKdFEf6YLX1sH4l
VpFQBabAhcsSKQ5hlvmzghjeueDGgWftu0zm9FR+6EcM6zh7E6M+OWrqNaTNYNU1UwyzWhAal+I7
h8PvVrWv6MSv1ibjqFg6BnlDAM3Vw97lw2qNURA/mbSymTdYlKiU4Q3xfslURb3e+n6MGzoJ9jCV
ps1ZyFpXdfFG0o/W58quPj7u2n7HwWfK93pzSuD07P9h4c6NQVXmnEl7aamKG6XdvQf62uF7px/X
n9DBd+qesIwawit2AGWE4aEpzJ3VjZlugN92e29Zo6a408B1Jvhz2T91pY8B6hf3ICE6yCMq+l8X
rvx5gsxQtZHHaQSxv8AZsGbeiv+mRP7vt73pqnDLMTFgQb9e8U7VkWQgpv1XQ1Jed0R1Ia7NL/Au
mib5SwwS3nJFbo3b+k3sOuPUPef0gHPYKXPuk7G+RF5OX3CQeKi65uDgqomVNO8fHoatApH9eadL
CbysTuKxkEkTpOqEZ0NuiNnTrWcbLFXDObY2NqLn2KD0p9Fpeda9cF3e6uxnNVfOAM3W9nqLXKCK
Amib2sjvJJPeORXGZD4FyTMPz8jpFSCf4+CnGY4JrwJZ++ss4haYpQEbKL7z4+1TIk91gICgOuDb
C+UOUWTX5pZmo17Hes7bq1sqfHHFazrwNdmdPHquatPy6ghJHE5skafbs/Al+q/7ZBGtRm2394hF
EBggNSqK8d2vhEIdK+w/h18TjpsQB3zeyZWeO+L8Bs2ucsbXJTPyB1EFWhAw2O65IZ7XL8Wm3Bit
HyHWi5bHX45xkSqYDVTS3bpkAK1BZ8GwUxIhnP+9b6KV1ffVIyu/pg20oomyzAHdY1r/+yEamahw
a5WtlINpCzH0hGs2kfuZy9VUIwfN+WbIrDQRXJDUbcqzcvww8R3MHxg1swga8oQJcSwyw4Bo5cJT
x0U3grbIGdsAJ5QIB3WEJUucZdS1KubLriNiJc98xmXYl/5AvF1LgEirbpGA8VxaDN+UVu8SUbKu
WLgJYsWNg9jrk9cRG0I1OoXfvVaIOXIXIvQIM1XRwLV3JZKDXo0Bl+D6zdbL5UO3zC7+9EeN5W7a
xLqFNa9trKFJ/DPqfYYFSI55SnllD8s+6I8hAyjNanS7P01oxRWP9K7LMlO0jdRSlbeadURLwhyu
ai9fcSFov3rxSbcEog/P8Fg9NtFxe42+vv5xNmRKWvmN4nN2NtBMctkHxa3XoF8yID+Cbzqek6YL
iJuNGhwP5LXq41K87aTz88nOmdbnzKUsk8dYSsj5nt2+aO1WIvT3NjRP0aK69OPMANCKQ4zDP09c
49uWVoZRwWEnJzS78fbsDxAd4layjl4Lg5Px49NrBd0+zjebODmGXwt9AEIolUc1dqI85CjypVmP
BZ4bqmkCzXZmbIrYKRVEnlA8riqC/7K6/81BYwpr2Uf5fDaeCDd26ETRz2zlzwxC3VXl/wrHL/3V
gW4vaCpHPsVFYjTA8/WuS6UkneSE0Bwv7NfEcu5mcuc6T64jTPoTrPJanJOpn7MGRv1aihVCVEeB
V8xkUw6XwKUuv5b18WSjJt0t83h3x/i99iRIuYw5AQJxDezvU1BaHa8/qcFOSI2Ah31s3IJegg5W
BjXtT39DFb6Xm78nnwsFlsZmo88DpAuDMvANhko4TvA2p50o7pEGWt+hNKRW7ULP9omJMw2ra6ZN
bPLO3zhI1t2mZg61TXdjdfGscNx0Q+eyqufcAM93gw6MRjregXxWF8LxnV6dnEjXlpbUh5RdelK3
YMBcZ5UDVky7nBu2P09/otH/+VYHIA7T0uAkRye8D/ICkCKXYil/40Kt1XV6FM4tqL6k033SJhM5
fXhOTDAKYasLdsZUhc5jZhapzy17MPnkst0s9GG4x86Z+c+dsEkmJ6D5lc0yH0+Qs3FNaAidmu+C
4dT0rOnYdZ6keqKAteRbU5r41vL1hDlZ88LZiEwDzG4lbGEL/Xm8Lfs+dWBJHTSHsuSEgEQamDXL
stL4Frjo2VzYE0f3IVNajtKS+cpSQJYpivfAQj6aKhNXSgU3t1JtVIj3ORzYJ7PnoAVrnrbuPxko
nHEiIIeIJbfz7bdF7xofveKTxJCmRIc/IrzZ/bA9OpvDdk2Oyw0s4QzguRBsaWpFkuigEVyktCKj
46GE1aD9CXnRAymN+vaz6WFiF/Xi5T60mn9kULrP6Yot4Is3O2C0odaWJ6hdkPz6QlRExSPHN7DQ
aen973HSo4PnLhH+k4pzI5dpnAT8n5IJBJjjBhrt9Z1l9uZVQh2BujsGsChIGNgplNOeEgvplHTn
zqqwnMXrMG2bOtkSLzpBuauBfx7cHLIcJj3jScfWsXGiedNk4+C69ZxEVwj5WzSmqR0FVxJ1htkD
xe2YUsDkNQOZUAEdYtVtfHOJsuxXC2ygBJRkxEjt+zPOlGsZyM9W8F4MTb/73hnxpjXP+X7ja5YB
E7WptEUwojLFIVAGNIVqlDly2f2ijX5rL0C/ZmfYUbQzCaItbkPGwNOyNUG8RcLd+o4RQCuFWDCp
0qHQPvmnIzAIYcAag9O+9b8lqtsk6Py5Ww51qm1gebGBOH3QcWcW9NopZrdmGR2jidm0MAOEVp1d
PWShDAOZyxbtgIY4e8mQhaaV+6eIp3M/vff5Ceu3wq65+0XZtesPZGYwFJZxH4ZjMB9w1dYwebMb
SF6vHBPdx5BZ1NizbJwioYqSPWMrG2jDiybs+V2zUWFnhMnLLDhd1jSIpasUNpKGcS9ynAS90vFd
CWWJqQaHQmxgcOr5oNkmJb655XtuovD3CwLSPPfzeUgG1zHqYZvzccBXoE3lkwZLq2ENy7h8A0Dr
fPWs2GvbR6Wcj+kFb6CSrBBNexNDQEqrNscilyduzSieH3IMjj4Nk3HY6AWpefBfV5thIUYM6rfw
YJ7iz3ncJ02nHOyU11YD51/M9vhOd/e+YDGkYfaSpjkHnriYOEfZ9DG+QCgBC+QvjxUNUqgyC0Fu
dk83DQ0UF62qotRNlyb0o2aS6M3AK94e5rpaffDOHmMHg0UkimZAx937QcWc5cZ0jeT7C28YTVFL
jydlhrSNvSIJoCd6a5djz/e1JWvefDKsvEbZFynFkEi7oN0WpsIkC0wctPWzvtXHboJaMIpsOwc6
qxfeSwRmySgqH7kwXbCD5yQRcA0inPNUGIb0vVe6IwdRh7lnd5UsA2WbpDMlptt3MyhaPyR80qs5
U+yuCKrhpCbKUMTqBqQW1bp3tx4r0erDK4+7nst9F9rYHu1xm8hsD+VB7DMcLuxLj44jffRcYKed
nhumEwOJscuIkQYT5+9sHVF+kw1q76BMplSSOGR1RIA18qf5f8xyi+qCngvqWe6Wfm7u+/lo+Wb2
7nVf/grDoiUTxEckdW128a1161aT7YdpoevoQ3+IZ7WmFVlxPhAZqV+pBZjTtJjE6T0PIXLYDAIB
C3fkYpoyjJAP5xKWFG1cjyKI9ssAAy6GofnwbmofkVbcI1Xjhx7MLvxaiJ1kqIxLhuw/v0PNqpXt
0IlDDIr78NLghPONM6POOgU1WWNfQvxqaoVixxp99u0m7WtolafP6y73rNO0qPq3uBn4+3CuGlbu
5DICjMXNXOoAi7eeDXy0xEy1NufIqq6Wjubzms6Tb3KNViiBhMt3OgYNQsrIEyUbX4Mg1JiBP7He
MMwvQKLFs6ZCPVpF3Tj1udzopqLYWvS85/bfD7fsldn5Zd3nlZ49l5to+Ce+AAUGNkNi3d1ClH0K
wLx2jkmcnjZnNxrQcqZafHHFtqdh7zgKHnccOcQJyhatvPeHG8VmxAjfE7TOnuLyoqAVZEecMgjP
t0c3kIlrwVLW81drA+ejj9qAiYf3rD6hoNAg7ILsWMg0crdAMrlxdLbsBH2QkIDP/3sR09hJRFjs
vhdFtCqDkDvxlT2+C3+ku2kCZnGuYv6pKK1AikFSvVxGy8NeWZr5W3zH3wCqUMMZtfWkqeCpPf0E
wLrH9UgKqBMjV04JhAPenEuAR5jhkJztJiSQ1JClfrEH5/BTVjnOd1Qd7AI6bck5sKnHhLw2yDZZ
LQ2Pa3Q9EOy1QVECB1FqO5ohD6Tf0o8W4TSQ/S7wMMB7wDFHp8ShotMepdtan32G84GenJ5hiKUp
Os9I/lP5/N9YbJW9bXx5LBj2X3toCo55+Jsh4haT8yAnUO9wzPOyMaw7SZSx2XNU3HBwaDtAHjWc
52Er+OuCNgHywwz38X9n0ABEOqn651LBYteJYlOhOLjpJbe9DYp01exNTloV6FkLHDVizuHkeO0j
NIn9c1rIxIfZeNqyRKwJc80hB90vG+14Qh/Fu8MCh6AcSDe+hsF1/VxXoeviaY8Uc16u0VKwEtmx
+E6VzJX0IXK1+F9Scvq3mPBYdUCL9vXmf/Y1wVsCQX2oOsBcoyNG/gWkf31ao3ciFKpXf52iWUsw
0BQmIR3OITkleWttLBR+uP8l303dES/urx0A6numQshgQWvCKI1dF8oacFUrAVN3+dnAuEVqxGgH
Ar1ZC/iiTWv+dYmkYHONuhekE68B1ZoV82XjcXveF7Iw4TRFgln3AUa5tnecRQWP7XiP/nrNN+VR
5GKqQv6qjGAu4oi3O1Y2tRsZUK9YemIBZ1+OJ0e4KzQkINLWfwtue2KCcsxTd6kphoMcvBZ6+wZw
hXncqkbdzrn0wrmddo8eMRjUJaYiIYHvOLuCUJHGyUcDMBa1+IBkDck4ullc7GZ3rxncumIM2FMj
H1QuH5HmXTfEjGiUYlX2+JchnqCbu5dcwRG3njiLi4RsJipv6yFlYkKyT/v5R4oO5xk3tV3dxC0/
MKIZgy64X/oTJQyXiRlI162Eb5d/xnBdC0KljNn851ZjdrQvYW8JsPhrfzPhZd6cAtDFK8ONfQtM
FI15P0ZVQK/CBPIIURG59PwCs1OjfOlU+OK+PFOQfhSJRFsW9vkuW+jodl0PuAb97MKi16QL3tH8
+KwnligLFqCtL8XK2KibEzbbjeTK3uuXfskTDyLVTvWwpQYIm4S+RnTMiEGW2gOf6cKft6JVr9ZA
1jj45MeZdVgjcEYo4q7T4TDF9QMRde+WdJkig9nJ+wwALQE0dtigt7SX1a5suhvQaTQn0plWo4iY
bXn0+woxu3rO97IELkXDkoDOFwyqVCX1UIkAkPEbvZ6sIjbhVujS1RWUznBhznISU2xB/Rm48sNo
2sRK57+J9vPG0HsJFoCPUNsyanzBXKCDRmysbDw6/ZMBJDwwKjlZwhFwzslyBAKddujeOZaIp9PX
PkyVf63UAJPsY5xsqOzXJYv1X+OvbS0Qod1ppuALtHjo2/21M1ZxNLf09y5E+Z73jKB5nLcPGwIY
tX5YyGai6qOw/YtqBcDsHtLkuq/idBjnhyU+Gkv72mzXLYFuBm3gP8dvxSLwLyDB23iLjLRJrR8l
wdiJs/dOiAm37sOAFaLvNypl/FrzBSZYlVWfq1xeyFpYZyguht4U6PXUPhAk/vu4xfhndqAowviG
sWfa/HPdk4LkpMTTB1Q4vrq+6wXamV9+AEh0sPnMpKfpPaWfgDWFdsWJjsXqO+aC82dTn1FC7lJf
IX5l60cf9DUi5YBsJw4iGdppHmQ1NkxYETnCJCweVMCDkiRBfrij8SO7ycGpoPBGB6qxWdZ9r2vL
/sSlkWpdpx4iwvuThG6zYyemp0/Ks7t5e/xNl2EMp4V0r6ysGo755RkGjudbxLUxflcdZBXiYmZX
zjMhCK0Mj0Kxko7Z1Gg+Slil5NWR/9nP0ffbmRzNQUOPzkb/37pET4n10/HgO8TnFlcO25Ose9q6
JccDno/ag8xQz4IcGkbCYUtyrT5c6bJr8dHZvLF8xOhZi7Z6a6dbyGp1GDCnf2hk5uiJVTiOvZE4
rmoJ21qkB8uPFbhgnrtgnaqx5Pq4yBraT0BuSjqbggCjvk6J9qOJBnnD0tH5t2jRdH2zeg/tSP0B
WpY7KOIgBuEOJBeYavviZjIU/vmveBH35g+N5xJrMZ0mRmuph0QIqBTtrfGp7/igNkzPc+ZgUHs7
k3AqqO4qTRh7EYRnbAoV6CoLBOTBRclM2qZ6JMelKi+WeIY/tckGDTaUtIQtLHY8PDEvh753Kmx5
RknNZUcukhr8Is1LLCqQbsdAOvMMZkPABBsn3raLG5raTx89LG3hSqcYh3qckbr1eFpGW97NTb5a
mJracQVzErPULKdqyGdc5RAjSzciTlEW1AGq9MHhOySk2QRnG1D8VKQKto9KSY8NRzSh7qCDpWIu
1npjKVThlm6NbfHrUbzGWYoDp1Y9kkqJQ7oy2dSbH5wGVEFu8Dyq/ghAoSpCB2yFNLtYKh4abNLh
xNdvhnmaacgD1mUruFQqJeSQqOGLpfnzNLs67gev4mwT4IkwGSxCT5lP9H/ureG8qNrqMT7F45FH
31BYoUv/S8bpW4NoJxNPQQJ0D4WcS7F8nplYfgLQt10RBLHktsE/6E/7jXs2cQR4riQu8dRCqP+0
qIL/icYGtdZ4fgvXJdSehYKAw4U5ATG68SMppRs40eMm3fhv0c9JIM7FueCjuRVJLGC2PWo8QfCg
swz3uhX/2kRbLbAQuM/tLgjincnbssmO6FqIC1DTkWxAgIVvaZT/F0Ydnsw1JrHmzWwizOBdOaAV
csgSyp+dAWRL9vOAjzN9GuS+oRXLSAWClGxmdCumPZ9L4vkoG4HQlXViH0DIhEZgEGA6flpAA7E9
UKQV3JItPS0hc03aIsLN7b/ZcjKODe81ikEvrXSQQIl10x1iSlIgpUy8uSt599cxNwEFkXwQLUKs
7kDXh7EQg5whjFVlrx+NB1PHu/lxPq57pLVluLrTN2FMN/rjyvbJFiXqV5HBFVE1SnM3QrCMpOi4
d7TJRseP221XzMlbbs/nJFUFvQh4XfJNrkFsoxw1wD/Qm7X4k9h7bD4X6QkWAf34ncsGvu6N82Tg
k+AgcuPMAM2c9m22n1wElb1GwyMIoAq67GXmTIe+NtPpZdcgyz+fj1EZGkRuP24Qiajl/opPKfJz
sA5K0UoCdLFlS4yqLiDW3MKbrfJUrQ6X4iWogtt4zFGF8+6z8B77xjE6CBPkMO70i8rwZK1AA5We
G3Ca7Vzr5579s2gqqV9OVKPXhmUL6p2aBQzsSSGCzqNLLagC6BNSQ0WQDkLAoI8ZIshcULeGaIQ0
FgVcRjoSgfbU42s0sx4p8q7iYKmdyPOwr/ubv4czQAlJfUn2mGowxeAwqDO67tdtJfjruMDtf3Y2
VNpxo4nZPY3ZorLRc3H24aF5qlvlTAFGrqIE+77t0GYKqwPRT4hxTrO0eH/RV0fFNaRPUopcQDIz
CmgXpIz3Fv1Lb1uEWYSGCCkCmAJlOLFK0jWszbbsud18dkZFDPcOL6zHiuit5ly4r1rpeO3QFj2U
DedbJuj7uHxakO+r7JkcB19HmOcaQ2oEwT2uN49Tg1bTE6sulXlXajMvPXNy1Qa77aMockjTxBY1
WW9CjeprqXXJ1uKJq5AIQyXy+yKTI6bXA4udg/ivxrvVAswZHKh1sXkl+9jyT2LQ0FJsLMZ3vbse
Ncn/04zB8A48KEv8jOHPuMidQ5BR4pvOlqszIbjbGkgT+Qk4dT1iDdC0ndtjQ35NETAgHu7TjOl1
tndozPwTaB40qIAvkD/jeAwqItkNlL+g7glIJ4MxRYBoTolmRuoJLjVTrGIDOtd7DbM+2y9+RDnG
Pdu67EURb4otHZI7Rqe4wpm8yhxG84V7mPyjWHJJbw6Uzv7JZFhm4CIbxbpmfgI6EU8AkuT87pgw
KAZakovphpCvhx7dXLdfsTE85bfXhplP2Dlh9kwm2ZHW6TPYPoIXCPsH0mz0cwYX8bRUoFmUEM4z
sJNX5yPGkNNUSIxACYqRcWafdi3aCmTCzhwEenZzm/uXplLL6CqI54Ci+ko93peQsYt3E6+rivFJ
PPMTsuctBYqxx5c/G1CsZBlGsmis95iKWdwCqrI1o0BemBgL0/svY7cIQXM9j2vaVaIeS1cuw8Wc
floXFNx0aW7RlxV4KfQaYL2pOkGuy4rJ3jqdO8HkFwU+GvXrXTzeQTp67m4CTNF/LgIcTIE2rWSg
NfG0U+rb34h9F8wDtUmk33G8/sJLdxNHXxNn5GFrA7U5GLOsZPjLjuOajXfu91IYJPjUpPp2+UgV
d8kuDBKvr/8s03b0YOjhilWALe5GH7tRvs6CaiZmRZ4OlUoJzAUniwsBzgb3zp3DfpoIVEGP0p1x
K6tx3EQ3FrpjJri90VcU1+LQU6mk80zn86hKYjOGQcsWPVCH+wP/aeQN0UzDw0+GjlPYELK40Xkv
qJwplZq2l01R2phKVEGelWKMCjGJ1kxvj9+N/1I7m3qBX2M3UB0hpzISIIlsYtEv00Uq1NiJA0IX
auAsevr/ETfWkJa68d0noOacSyDGNZaUohpnsahcDYLy7B2j9O/YGU+tzcj3BuGzppX8yiddo9bQ
icPhq86gIonDcfIJK6lr8S4/Dzn3zmrrEy5ZDawHBi9wptlW4gTU2W7M2lwD+cGWtP9Ua4VYWntd
kFXt86fYpSwCxy9HzP8A7SzCDq+Cex1ryJ5P5YLIplqVgZ1sJ7BUPErncJQoO/t6phuhLziolTZP
ez1ZaWQUQ/T22S78WFPDeT3hJ4WZvbOTFX9Y6cEvZl7Igaq2MRkvPk4v4ruru31+hzENxcQUHsTz
ZMXtzGYPKcqVqWF8e+JNv/bbowPcu/5VXUNCrDm4IZ97c1JllaEW7x3lMnSaPBCcniy2/V2KLZmk
8fTEO6WwCIBIA02pG12tLhkLUp+7F0FE0y+mpmcRpzhMpk9Pj5Qs5LxJE/hESTKltZ4FAgnMDsmO
UoODaIxCLx2xFZWRv5GsMsBKEKBqW8XctjdkwN55P35xu8kFsYEoZg5cAqdDjZEY4VChRvQu/N5i
lCeO0ZabhnJKf7lpDPBAoMZSjrkHUHyLqZGPhHaXGnWi+ANpijfF80/3bETkDFtB/kwikQLiQGdU
OBqu1ZbEUICZnrpiphrC1TEmeHjz+XELxveuub+5G0cMCMGvvIpfznIRP/6tWNlMEzKgpXapnxGn
4nQKIsx4atuVU3lL8IEF3BuXvtisI8zOG46PElHIUiKp7QLKverrLoV2ZeGMVFNixLuHCy2A75ky
Re1JQvEAf6Sde63IR+oIcfx+o9KapSUHdsRFNbubs3jbKElyaMKQeED2n0GBNpTMPwy6bd4g+KSn
yWAQ9Ts0pguOndu+h/G6OfFkb11aEF5cxY0eGpTd5IxIhJP5fGtenkN5lJWbyzdGwuXYOReUskVE
gIJmo4x6aUt/vX84UIwy1PV6WIqRVA06ROxTe/hVY1oBieTp6lJqTN1LsWPOgPABpQoAT0h9xVyk
OX/26j/qybjEjEuZSxaLDktamLQyN3idLgHv5UFOoZJv/MmiEQ/Sc1+skJrFVC3qZ4RAoEOrNYdG
JdAm1bLfVC0HCzlUJSQZtaWt+gwctwLvGZqva4QQQpREPYaON8K5N92uzw+uNglVI6qLEo1vVjYA
5qWrDgMT3pvNY/nvczGTVa1RLZwmn08rbiIiO7w5szxppr20atAquxIFMQJU1ft0+Fm5BweyfVAn
V3bNarGdG0POvzCHQFLiCt+I6NT0yBksvMDQER4HRbt4Cg6isrvHNKmZPi9gkEWC4mPxo2fsJzLV
cAPkHiJKMYB4gX61YC6tx+Fbe2pLrAR2z4LVcpEnRAn3N+XOnLTpCkrlTZ7v57Z6/XwWQdUpHUpB
sWgB7f2r3S7VSKKF5a4Mc31uaLYhzSEpLpq5YtvcWY3X+b3yIik22K173TdPhOlLy8X5Bj9wgK11
Y7mn70KDQv/5S8ToZgC6sQWqg94jqg550h48TK2MNe2F/ShxJI+5CdyankC2FZrHWiIj3gKvFRfP
u9Ac50wxBeTAo8WEN9AUoQexXyBf1hpyX8ztUOsBLU37xsw/yIdlz6wpXvpbQkYLFkpVcABA/fio
iT25tULu3rV0vLIFuwvDLvia3Rbui/TE6KAPSP+FxOdXP5bFDnkqTBp9JDGl9oNitFu4L3vKDFce
nSOMZa56xznWTbsLfLGH2zghzYy9n+5r+m7VZ3g6hbpAmg2IR/xeQnJHlUR44i35b7Me/N3KJJsT
MXg6TrR9r5pLfWvYcpVdHX3ja6cVUmg0kS/vws9TPClDroH1hCsl/lSKlnAzns2dcoxbxkX3BZjC
H4jSfRrG/gWUXu04Rs8JrMTR3lP2ZNLJbV9XykM4o9WoSzgJfHCAbtKamBmMKCnS3SS2Ftgd71qc
13Quva0Ecm0FV/OfE9qF2giBYzlc8fb5MfLBIc4adXil684+U0ve/FK5gqQLbV0vL7KnymInxHj3
UVMjg84KE+GR+GkZPaUG62f2POVEy26QbjB9p+ywrPQZ1BH5mTg7XzYtR+MU+KOoLm2cvqL8S1qO
1aagUgJ4X15MTv3EwVsIE+hk0GmvHawsHX20qN0Ncu6EqC+F/thipp615M+PBPP13WiR5R5Wz2Bk
RaXkPSwuL9u4f6TTSTqDSBowXd22k86glPc3FfVyH1LPUGIeplfWW8Ey04pz7FguxJSzPLQThxjV
gk8zqqLgX1L7l5W4q9/KVM/ov4lFXO2Wri4J/xebrAwqV+91Hcu4Q+yt+nFFP1xmlQ674yet6bf1
nLxqNp9OBjxypbhxp97pXTFyOD/INHo1J1I4qE/3wmuinyHI1qwVsSh4eUit8r9h59ZyCZ1FIvqh
Gl5fN7Cj77w5h3brPYITA3sWFLnUs6hmxEUd5bLDcwsNGtULCsJTjqptSdlYC/+d30PvFC+Lmy29
O7SdBe9S7KYTSoVQLpUw8/zemfWCono3Btfe0UT9inewatleMH35a/fstYxbNsRrh1fqLX9+JG3Z
1XCtyEEtocb+zKx7nP66uA8Rw7jJmuGrHL12VABRApFU+vTbFArf1esgNqO+tvw09ePR0sFU3Ytv
V8gYMRgK9t87j81vtQD6wZk5GcgCW9ca5m5RJB5d7JSgZVd8ngedFL9b/Op15prZJSWNaUDk147K
85J5ZpN+eEHuDIx/WAsnCFbcwsEestNLpGV2yo49wltHcWpafhvnRD/2bWTxBbmlz4EPdCMhqUBm
FKzNBPoLpeV9On3tcvEORSUakCURVr138S9bYNfT4Gxdp7Salup6a+1pMb98z7gNFB/iiPcZnP47
xa6P8GmUwt5iik3daDStcqxPLPS6EkyW6U5m3UpJ3qeiPSNr/3+puO7BfCk1wbjIYARHX+x8m193
uHNG2rMTlXzo1CVxwv7OxS2Zkq77b5fuMbX4hXqaz6dGuubwrr3yvUnKqCSyVeuVMtrVeCDHoZeF
79tVYP34VYijUo6/TeJy4tIH9g7c1Afj09/wUa99d8P4S5ZmdW2Y7NqXl2ZMKJnVnuIOODRl/wjE
I3PKHnUjCIvCX5PhwGKZxUOLNc+opsIxCX/6ILXaGIXKF7IfZhvU/8IM8oDk40l59afWdUFkpu0v
sj4YA4K59BnaYxRS7TRSotH/vUDkE2yKIBrV9S6oPdIcsoJfvT3pQATjQ50eacfefEK2MXyZoeJP
LrJuzQ7PrJak4esiEKNNWrkap3J4XdPORK+9yC+RtP5LKTo4MnWzkoOCapOP+5v13AwC6ryqkpeb
f4ucdhGsVAVgQkmQEoNpZaHhT77WdHSSsizFQWnRtleGMBAHiFWtsyr1SW5XBHZjT3LyF/tkqGj+
ZXNdcaRQVSNZxZxmYcABx6O5o9GPJfZOAGMLvG8VS0W30iN0c5iZcsAZcIyXSAyB5xB3uAOznKHh
yIermoshWx91mq7Qk6EBHs1YynWNrssjhBJqK8nYM16t0YTFyMVi4hYyu0P9OpgEHzEPpdOCkBLc
MVwGr0/Hyq9zmhRSrp0JV8MiCuJm2AmplBSkp3YD+TShQSW9L+u6Fl3BKCpuE6XopQRB+4ijWECO
2NIaarjziC3DES0/tgLfYpmuNBankPComxQqeHpta/KEymbXCHPy9Im8A1AojGmJpZSz9Y4w2s9A
Q/m5tTxQh08JrEA+a2Ai/8/2ppBmuW5t5JMv+4oK+MnDOTTYckXk2KCq7bvb+8frACNfksTRpgak
kVi9Sh0mjcge3AxCmCck9hwnByWJQRMzzitMRV8iIFdhY/8SNYpfq5hBpfk2coF+Axf3wFKJEx7U
KGVv8p5+HlRj/n3MTkY+8zdbHE0v/5MrTt/1tvuENwZ3cTaw9xh2bLKWm7gRVnHyLjfWOIFIA3BB
aS0Vz37Yt9LRrO/0WiJAUg69sIahkDL1i3hD97SKcntDWqC8AlYVYRZMoEwSqr89BRg03PY420qQ
yfJGA/Dp71EnKxCEmzTCiuKLmmaoNpd+pT6AIS9GP0msRpr/FjNA0wvwGRVDJp0vBgRaO1v4O9rF
9R/6IouUg7j2kzvXvevFf6SCvECaHvcmaEKZutAkPsjr2Q4ihztP4sqwpC4ujbhB8M+XMxte4dY2
atg/JZgTSAAv7VN5F8C1YX1ltre17qigPUgJK6dP4ETauTFjHFlh6Sahl/y26qH8jQj2mVkKzRfO
ZwAT2Ohx6iCQs3Z1ZpBMKIH9Yo+VacWT1e3vkn4CKbyC7e82SXc16CW1HAJLXK+H2EaZ4Qna16D0
0vU9SF2vk/hkHAfi3fPa+5EiHL2bfvcOqyJcfscOtS3zcDnsC7L7PcAVtm26Dr8VSngovCBsixXP
oneITh6Cd0UWGTf3eKgUGqcsmbHAfdA6SbmNq7kbI2IN6H/MB/Ytg/ocroF2sB81ehgbdAHaIVj7
CROy25qyYUFXApWGvIxZmmZnpp/YFFIxUfvzW2cYPZXhq2vYEg06E4sgIIq/fNJ4ZpZJPKipIT57
ARrgJogtZTpD9/khRXaxpWwGjMWEi0XdUoaSifUpXeeZTsCFV6cBbbD+ZZ96fPv0D0bMWbTex56f
1eJMIWY/KNQAsrYeqJ5l2KmHOP5s/0c8YjfUwBagv4ynG3nfp8hWUriSOBWQ4DPVXJD5LwsxBXQg
8fPb4Pf6Dicbmy+KKZwQVjy714yTN4KOrAKC1uAiLsI3iT7MHh6s5CCxfxRaqx4XcU45wb15QWtB
HGdTl1QbUGInEM6a04T0lyToRrWZZ4ZcxAOTVk9gvS7v7NYrbawffR7BjKNalDBIqTurdU0hD02m
Tnb1XqKJFHFIYX4jzT3R5Dz+xE1aGk34cd9NXFIq07bFsBiHMGScKiwma2nLpV2y2AQfgdw+cTeA
8sW5xcpcw/qO2rrLcRUAOtJKBY52ls6hnN4mcujlVW4IIirKfICPCpfVWduElMcdTQZD3pWvFtUb
hPUN+S6Xk8MLsvfket65ky5c2Z2PG8vu9M8xMzVaEz27iN386e1s2LssfI319gT74YdCUGKkNag+
zZwjpTNeq0VaOngklVUdHzX5V4IVmGG9vr0vrGSFIZzRaNkEJALmWCicPDQNKjVaetpGEcQe32Oy
Y+xgWQ3wsNUc2ygoC+h6hQEXcCuEYajh90RP79bTi+wZt0py73h2JjH7zcd2B8rtmxf8unX36lLd
ZACAhFhUzDr6jlPd0TO2v0FPaEbB2HvUc2MLPSeZSp7oWp037qZU/+1H3najmGOxvQs5ayMZBqDE
Q7/NmLHk9ZtmhFlkhy1XXgwDlHlHqwL3OrhcGuZzOD96xhEJ/WopgGcxz0xsZNu0wC+7A+ZrzTnr
d+UHg7/22vmi4x3beCS7gwwnEtcY8L9rxCvyXF3wQxfrD03qv8Y2NUZfHoredvuEesvRiSI1GkMj
UzWZRTLAJvj6xhLLY6YkEwZMnRnLXAJzfg1GDyLCvzDklXWfPPBfExO6TzUm4MsUTcIej+oKrHMR
xXSElkQ/I1UgDFEk/C5nQvG7p9T4mh/fZ6BGN/5SZrnPFyeexdmzJJIGYNlQGm9X9/w2mh9SEQWe
SWr0QuQOfcahI9xhg9+rHYGk25EEYGj7GDvPVqi3TcAJ6WSRRz/GVYddJMmvRUgDJb2NHbWbct4/
5zI9wOa7Q/vjq5BcBNMomJ8bF3HN2mgcDHoA+i8loKnvgd7PVQ2zuwpGoadkx2usi0UWWAZwY9U1
4jkktOcvP6zF+kQKxDmpcbgG+hnuv1fKE08cc7CucCyAgTB8Jmy6IKz/Mfk4/h2KpPT/3pJkAJEW
ROYEfw4/2tvJFm8j0lsbAVob7eFY6Z6QDne0meEilDs0J1gAr8QGR9StDEAVTOyD/zRcuXjqaP6n
fi+n5Fpxfmtt1q886LCAVGiv+//6ShPlQaa8WeMUXvo9HLqnn2BBcnBr2Df3ZvsEG+yovUXeJn+8
gMjooqxlExTsUEeHUYrUWjZMDHlTyhQkWHKcPVoCy5t4pPwEaTT9iHedlhUKX/R+ms+B6XZycqbC
fa3ImgOcuDserxh3PeV+0fCJW46zdvN2ESot4drVoJUm8e3IciW0qZ3byHexNJs/6D5EqLtPMhIa
BttgQhWvURN2UQ5V88fBcOPmNQg5tQ70KUB5V5H8ljF1hwnoYjL2LV5l36IKO+ThwaC305U+QwYU
GYbgcjlyQB1xKu0ko/GmDIRMuI39d4RZkQqJmoRbTxvU+jWMhOzcgnYo+RDZUjwR4am1SGovOo2v
iN0Kq41oK1AL3PjUpYuipht5RGLsq5ON2X4kuHE+nibUkNE6hqQbsoBH7UJRThl+j+bX5h0K8bRp
52hqzFhoezxbOmvOS1Uq4uhXQzQKk2eNaHhlgsIOs69JRkJY7WH/OxyEpnXukF67rSJ5/quI1rrY
1RCje3J0o/7bU6ovtqTwnOojeigPiV46LwCtfCblcegOwTx9m2zQsqXsaMvJYAtP7POdnpEG3wqd
AI99Z+/1GGfn0pcxJXA44/AAsqfFDNQVE2jAwa77rm0MyjGG2yp7o04ghAcA62zVwIgNKFbwYiNl
qvm0D7/E3ymr+HNpWn8PwPPn47BZgcyctqMZH1cBUF2Ta1hCDTdMACJYPUl/47RtGDVU8vNfClJA
Mro/Jl0sgiMoWY6Nn5/FLAceg6sEWYbGrsSd0nrGT31ps6nUFIc/xhAsWvXI8Vv+0U87UNNhQLpQ
vJjCW6R00b9rjFEI6z5wx2+PuHtKhLxN0ZP19RJfg871EOsIQAaOfWdfesB9CUrV7IOAex0Z89ZF
ReNOLoIPvRqRXvY45GlcRQwc86apTsNZyy5GHHt4ug2/v7lIitSL39SryAKJgBiFqsCkR0JLuJub
fimq6vc0QLxmdXFLwTrppyVIiIaQUKGRL50h98oCDVgHyq0QqHCJSdsp4+J5o0JKK2Bnmp9Zirqn
gVaxz3nYrTtDSvaYC4Zgvyc9QJDNz0G4HRyHfE7S1NjcdpHnoe8DzXof0j7H+u+AsK36P1890lCg
WvGRqjcM9Clv1jGCau1sGISw3/vMMOCOr61ntDLpjrg+DQjzs6aJiLSfjgH3Jb2P08YEbBDfo5eB
sanWPFXPwwK4wqBWy42OiIZPe+1z5wry9ecd/h5g64T2/HLLWsS42qZvdxw1FHmVF0/r6N1VF3DE
W/vi8dwHRNKxeApLjnV6VDWHgErEaIijWsoTGaqJLEbNSc0PCPNCfeGWlhzwYRPRcb5xEZ4n54R7
i5jIeuntRFuJEWl2mJHXei/X5gOxMQZCVAMtvXxv0kSkSoZ8c7yHy0oG8OX5kcOQNXV6ZrZCNcAA
r1sy79Ie/tGWUEDLG4JTi0xBnV27rAOnnHnm0phvqN696bv91rSPYZ5gIpw9ql6g66EPQ5VE4by1
fYGXtbMb5tGImZMwsDzHxF8N6gEZQCnsJaqKgR3SuoIgZNGL0HM0/ykeQ6Sr05trjROA43p5IP03
G/4ChTy5e4Rc0sz2BkjF2gSDVMqLiygkXaBOIfiAbHase3k1tDR0M1OiEeAKqZvjfcRKnB0P6p4P
zQz0/FJpRt+m4KLMRhNaojp+Mg5SpjhNdUGVUGa7FQ5y8gzF1D+RyTkWyAi++Yx8W0Qqsqu+ywOv
EIUdhGH5vy7PzmzLicTcAjsSVxUSAh+qXsx1zCCImuWMtlTKvCqXV9P3O5g1IOLxka+iLWtYFBsj
8ybV6nd3OTxLBaJopfoo3Ychot4dXSRnCrOWUcDv7YHuT6FLehpqPU6HNqdiccdVxZw1h91JuLn+
ifLv/9Y33OMdBcBBhlGum4EWTkbligBygbUaYMyYb5+ymkm76MJJsbfEWy+hVMBb3YP5FTvHNIoW
7/rXsMXI0uy6JcLhMfCYrnT5CWomqGT77KCOTfaW88XoE/yYhodBx1C/LOEHNz2djmMsdhU4MsKW
6NT5FDuTdHj1PHkm3YO7bWaazqp2HH5Yif/23SPpSTxpaOAU/zYccdBt9uUMHldP2qOMUFTj8jjk
rVLVqTBFZTln38s02bqzBMpSxZQafUhpe4jRVUmCugoWKKBDpQU2CzVPzNGlz9ITogTgAHtSJVrA
o3p/0EWW1gmqfL3PkysjwcvihgBYO2iymX/wd7s9R9xdr8okGvyKM3giLFtwbgj3ggur0yJOn3BX
HKTyWTt/OrXkRaqZQtzpz7At7mVzsJxz7YLoVSZr0bwftzrjV/piPO131BpMncpZVEqQD9YvoVPh
Js6gwbqKd+iGWTr3lGVsfGzXG20dXtsMKG6Ah92b7NfcEW4m/J03yWn7Bx0fozNUwsPP5Qi+qLLz
ZXlmfnIC/ijLWAMDM321gAIiyp2v2jhOFwrTIke0usCdLw2VN5zHwguDjBVbkKTNUxSRu1O0s0yJ
P6Hejf87vDvGqVAlE/ktkP1oHanlMVEou/3FK9qYeRSM8sIiqUNMY6OxedtIZuoQQ2y8mRUwjaML
fPU/L9WsBgbeg+VdgYbUd12sPLNZ6rhNtgda4FD6y5GAiGgSQcCwxzbKUebJ7mdmrW/Hnnf8ryP7
rq4qIXjSgss38yTR1m1XMmOodCQoXvOrxVV0WfAhF8T70Guv0HAYiVI8BLLOkZElolzMa+leTBLS
LHGQV1/sT6wp6RCSDgvISLmuI/xhGg2dOXVQBaqSVq+RpTeL+NlaFihNCfXLUh5UxaHwgxsPoGpt
w6v5vLQbtNRntpI9a/tD4OJJds4NN0NRKv7lgGMXFQGj+7ZTiaeBlEvafi3LGQRwWBbJOGYx2Uck
adKVBZz0Anycq2J5u1ureAYSB0jnPDwHoTDwy8ZfYThCnizsvTqc1O+lOdjroNw2ZvjkWWCp9cwH
DiG258ugu4EIk2qrcgXaiNusUXj4ezmtTndj2o/8e5kmVvHBMzRZytnXCkPZZa5XzDAPNugvSOSN
N+RrCDRb/+yEv9d1rEgR+m/ayoBMTXTgOfnNAdqwJdACw7FalTY0SrHSJ4dPmiOhnUeboTMC6Ag9
yJ1GMnej/q8RAGpr/5laPNO29QXg7BZFXok0otqEEKeazT3T7gu3qFoLJIxJjqJNGKem0gfA2m3w
00TR6BslMfzBRHoz/DKATlg0F/CXXOhz1Hk19bCm90gx9TMGXKem2JbQjg2dMVgK4vMbkEqE1SQc
f3elcsdw0mNajDqKh7qTwSfRVQ3COsszoxABmZf5Rym7mWMQpcvBrVyLtU8vOx2Qkx5yM3D1bqxK
qVK/IwiSHqZqRwWLvsP4Xs82eNIy0VnXkeFN47IgM7n1zhQ9yGhz0JPiGzRuYkRSdZglSkKArRkl
prmshMGAQkDThCJVd3AkDbUz4wAXIqn6kInRO6blm3lXsqhWuzjbXFiRIy7L2q5goIp3qT2BDMPz
OBkhoqAoy2u3oxJh9Lucfki7S622cakn1MFenFoDv5kbWlfyhTeVkuP2B8CDDyxhuYIRh/A65vxo
5/MgfGjFJkHY3/Bmg1A98rpKz1zkMQ5BTLEvkn8D4pnnagneielhnsOeFevd4FXqA5Z34lyrDuvr
7iptz2bnaJcGy/HFMQ+R6cp4hqTEpAqneI+1hrzV3wWrZL7cl6GGnNiCEPITBtXaQggkCpmizmZY
+Apc5FlsT7y80eqnIov51qJL2F5q7M6YGvJ5yeKioBa8+VgWVQQGV1oGhBpUcpO689C4VaATpRIQ
Eznee+ipLSXHrHjxOrgNT6vPAgszWnrsm8SmqmyQmTooAlGdKjgaj9e/T5p9V2vFfAFSoLO13ljT
nOTIqNUyRIz9SvWI/p7KVGnB2kBjBQLO8n6zwuZ8vAStEWv7XUrltxW2kzDO0L8OIP4TtLXPMtIb
6THh/XvwCb+1MoBEYTSqf/LFyQ0JUWJc48nv1exLISC/MRKc9nC6VmVUsfhPrizxlm4o07+mH4iJ
MAWwLCOHK7rDVZLqGu0X0WbvDMmC+Wuup/SVF0f9y9lBSn8k6sCppIqQJWmym8CPZf5leqpfOe0w
sQvCC7R6nxWfB73ClNnj1V01k45cqBQmQs7/QC95lDV96mns6WqK8LeG0CmntZ5T7W89TWCs+9/V
SnDGmvS7EuekV/R9YF2lZcjr79zNIUljGmzrHtHksUg5QwmEf3nQhMjTnb8C0S7RVOquxZN4AwTi
ziU1b9tCd0bBpLAllDniDyl7NU4fXQL834K/vFl9UcN1ArY8FyEFi6bjZMbRzVm9FGKHvt+oJiHy
G5UHXRREUxj2BhA8HG1GYtyWWIRA6ulZFEbO6a5VSbcKIBeKEMzRuaPZkuIWwkDmPWRxLbLoTe4e
tuz4DzXHz6EYRt/UTfvzAPUF3MkZyefKptF9ZhbPqRaUDHafQKI82f31q+oYe+gBGm1fjwmk9ow6
49YDG48p3J1zr6C0oiULbHCa3/YJYOfHI3wKsKmvVVUw/Dqsz1zRKRS0k0YiruoJRM8b+zOdRyhN
IeynuCWixXhoQw1BlZlEqkgLARu+5rnXseNJxXHi26meo43WMQocjuDIXAVajF6qi1OPxB33g65k
p4iOFFqsPti4XUNzh9OzPQsXbU+67EQBcytZWkn0RqzQ+Ay7LrBV+j9xZYsieG+pEcWNhF2lgx1F
RLPmtW7YMXrn21/ZRJp/cbzQ04AI/6JInH2jiDYHoGlaV1+dpTPlK9uBmTSoS2I2Iexozi8xtWCH
vX5QKiS6rnWHGXqgj/T7Sopqi7YL/CCEchHVTi1g2vjYexS+szbDp6/nAuAhDS7B316dMpqDUJ7B
ayCOaSDS25zuVfmVbXk4IFlyu7d57TdaxSYyXT5Zu7o6Mw8O3UWqrUjOFGvXixUPb4m4uN2GoWxv
ugfx2Jg5mP093nrlLnBE3YHlU5d7sTefcGG8rIPc2DLB0fltXXUSoc6C/sf1R+on5E9bVuQJzgv7
Ph2q5imdsHSfvujFcFS7jKrzAmiKbZqKUEzOndU6k+VXyTBGVaM8klGGIIM0lIEGH6XIJAmLWhFR
rkIDD55KFrAHSfQYAvGZdmfvScIZ+OX9RzRTN3MVIWpI5oFBOGkOJo3OqnbF3ULCcQaOtn0K/C8o
5irLWngExOWO8BTvBwg7uUHuX+NJNi4KjfPShQEVMaQoCZ8n/o0KU8rLfym/pFz0hnv1rmsARwwO
2irZ4/jiUrjLZ8DisUiiNaig6110iJsR0JDiiPhdkVJAPizFzCGBb9BEdy7ukmPx3X53AYMS+ApL
t7aLgz++fvH0guMurDtgy49n98DrPE4PdphnWMyIJEnj0OJ2OB7e6Jy02UDTvqzLgalJ7gtB3uUN
rka3QxmZCEJ07UYXkLLfpYPPAEyMg0FgdAQj2EWvN1Seo8c15Qb+ZWUk5QpC5qrR1VPKoQUJrJ6m
59mbccX4ZLGCZwIY/bQYCag61tFmXAmXGZTPglbH0UJ1F0Uiqrrj8u3bchuVwJueZLQlECIcBzxT
8svc1FK+b9B/obh5iIiDnjK0uYjxi2siXi/b3Sw/wt3HUk9j+MPW2blPdxX2Hvx0VfHDPNv/xQoe
NDfTpyAYb0HXJ24JON2oU1fKFZOEfbqJ35zIQJK7vLxoHWrY92Siq4y3hhe82+bBeTvECpcJqtp3
EOGUH7n3sOQzVSISmfUTxm70lD0LtiP0BeH7hgTzx8lRMIOYFF7kfWLY25RUo5eo8p/CxX2abZEB
OlyWiQrHPlXFUtKdCtzX0+6sJJ54PFQrcAAeJw1Zo4liel8zPGnc+kbVn9X27Yo6iCglxINg9daj
6bRSM0lZynvnPQ/HrmTS6jI45owRMNM7ohIB+Jz/kt12XmQzb0LYsjo6/+Yp/5KtiHBLvV4NHbUp
KUTA8btKt33PqiJt/MDFS2p5bLr2qjvJHOqGeJUx2nOfj95JtGrYVG7/gGETl0UFDc9a3n+hjuSG
abKBm4kVRMedmRtYZyy5yXTSMYgnqpAzfn64baA4ARfIJsxNHogVtCojHBqIdbyMns11nPsOr0tc
h6t+n5lp0jdmWEOR7CflprQ+eMTz6+LMQsbkU8AZDMViXSD2p5p71VGFD2A1rkRafvgDZkV+v+Wb
2IC5EcEEcQWy/iVbIfirqXWpkBFfHOMalnhsloA0P8yhND6jK7TVjEzoPQyk6hLzhz3ZQ2HoweFB
JfjYCowyqpEL5E8HRVManXsolCNf4AUpGuAiv30MxRd+oUjlbuzAUG8LPIj9yuVkHYyzxRmSu4Cu
bbZZMTStTpSSUConb64IME1El9TbtnNo42C2BNwLCaCYuUnqSIbfxC3ELhljteIzIHT7gR9kEzRU
G1Nm/jWV+MPj9GyQu1B+R0faMxOhj0lUMspgeU+OtxWdcRFpv5ZXqxbDf99yrqAm3Jxz8SKzNAA4
1j5c2tQScgHCKBumcysyG5WhudUy7xVXGtiBzpSI0xyDyQAScCuyzzTucsa2APNSRqlaUCczFJAU
nJ0pBU8YRI3totN9v3nEuDP0gjX2wcnp0mtuy5tcfQWVCMaoC/ZaobRcd7VHBgAWY/Q0E5W4jnyf
bwbLaKOLQpKz3dVdww2LsdaVLoDc2zsKkA24kNmI2uJOj8Bt86PUe3d9+cWrBrue6DnJeUTrKDwC
H6hLYGLu7P+0f4P0R8ROUSAIIKbmcENTti3VUpdAMLIdgX21AetQeW/yNX+fhLuPCfqgHRm9tVMs
IRuqBDYEGGTNUo35fjYkkC6unmaMHQfAQi/Yw5p/g/DFua23MlQjaEQ43F+sjy3PYTc+NmFkcUqd
2iV8CC/GrIqYPmBiZkogZ9mXHn8a+SsPW6hyT/9McHQWSBrbFgce8iLyEeUNPWRcxFoYAKanTEZE
j8ke/Xt4GiciqRNLUCKXH1Rt+yVrLHCrz929nKkAg+C2kuyA3Q6uxd9JW0GkICau9dExVUnMNedA
PUSHrrF3uhCoeiCD9Wy48bWsdhekRzhrkrkRmB7WaE9VgvgcDN1SdMclE371s90G8VWRqhkA/XB5
6T+D6dkm8uElvoFUGxPt0Psnx7Y6JgqbA4zEE8pDPnBxQHrkL8hBVLtPgJDZQbhu7NTyXNjVgZ6W
NRCWAFEcolbFxEUtJiGqhKBI3AzEpnNlUOPjOTjC+gcFfUgOjA5y6J/zIefW4yVoiXG70OXZjD9N
U3Cm7yn7HjJaINSZKL+8ultqAmIczn2FVTs33zrd1f+Pc9hyAjGGEATzMGn0Pf/1nJFQljoGY/NB
4uga7at83VcKDzIq5h6eZoEn378rx5onF3cZ2ovZrHQmpBApumALd5fQIKqLN0yUzJNYHbl9RBhw
cQF9BI0DwuGejvhOLypYnO86WVRvRrXmJDCMxrlDVwC5J0ogRCTWZNM5mAiD8XJ/aVmjpZAVOjFD
xPHcKTf4gCWHRePwrNkPZSPB4HzL/CoB7qQJ7acI+YXjPG0PodLg64dZn27mq2dsG2h+zZbCu9Lo
fSZ5HygKhAt6N1z+Ltrz4RVOAathFAFEQcTBwriBy/JFcjT/+my2/H82G/PrpU3ajXlRdHuuIqfo
E9eoMQ7FvRFRW/lXSdPX+/g3xLko+qTlJpifAqAN4bKRi3tTyyrd2LG3WOzbosGb6FAZRrUU6q7J
/ZZwCubAGw5sAgvI/yYJR7X9NExpcUVVOB8Grsa9f/FrSbwsO5UzLrSKLj3fs6Pw4oNpuQZjxjOh
Em9zWMDdKzB1mUhPDsI2+wNYc1NTaOnVi5doPdAg1DMl14n5fXNH62wLKahG+prykjr+Rjc0ZbSP
qOqd/qX9HD7LIAxm6DoSUkxNqftIr0C8QeGNYhdTCWOf8bEONQVjJohF2KujLDvy3i0ldYzIPEsB
bMR5max4jHnVndRQpihk5u2zcNX4sTqwR5kJ2i3zhMRX6pABQmJEN4Ado/wey/nAvizMlrMJL4uC
KxRBIn3rTiOEFePevxKc0aW3JN+pWJmr79kvCFJeE+SMDUxKJVu4wjJH41dJuCKHAAJGjGEHdnHU
puvzO2nANyA9ogoKZCNjxoaf3GVoIGnP2wbCkjgoye0BOXgi56MGYqwRe0Y8cEVSfJ0NWIzpcN0O
1HnIr6w3QJ3MbvcT/g2J+41hOaUOYkhl6C83s3Hbr1M4sncVdajZLl70TEWrIJsqNuuB8A+63/ZD
FNrmfJeQFlSUWASicxpBJ5IHdEVYcU7FKZ4tRFm/mhCLwGFcJaCdVPNUbJrihdW5HBtLXH2yDdDz
AZFMAJOTM4e9lx0gvrw/HwtvyN2D7s4ruHAwh3dzq38KK6kcbbg70+80NdfFS1o9ZV1ZYHKLJCVM
SQGD3Uz8sP59CzbcOtzo8XfhiG4cbdRRTLVU/oggO7e8RRsGASyHhj63oqsH8SW5Q0L7lG92hQ8y
mwFT0ago/lNsfCw3VVTZvqsQvsHOK5voUBR9wLy67nCPnf/TM7qMJoKpcmMPfR1dw7r9TMfi4TK+
HujdrPb5Wp/0JtZT1seXYCXhpsDgimJ2XI9ZL2aYA4EpkV9LSUmLU2LC7JN8oWOMhJ6lyz2uqtCu
yIRPs50yTynkZWADK/tqK2JwDUqasjp8SOFjByFUPGJG2z4HdnYvX1No6tB7yD4U2J2er5cUzmHo
atTZ7421EJRNsgh9YL2VKEy+IvnEhzgWBKvtKe6hL8gOLcVIvZmemvqTrYQvDQu51Iugq3y7TU40
ZDvnNRxh33mX6T+eY03B+poORUjANUxs24CuhKi/PbxtXqqZ7K0ObCbUI+7lP2oOGde1i2eNALyz
wr0H7OgEDbD5HAfsxIHO/Eu5YNoyQmHrcX5vJR7Q25MfX0mre3Z1KKVceuu9fJaVMyIIlq8JqBnq
ckCmM36nK6gInzz1LbYlyUqobX8g6z3ELAeSYjl4Z9mH9stA6k5FWXbvMpBO5eJKmXpiSlumC/PR
YLHnjoQdtd18vA82vdNvup8SWpCa+XVRcGqWhJLge2g/+CCVKt5YuLhaEEecsL0wZ3y7+BTLsQCT
dpYCRaOxOsyFSSY6qH76cLyKXJTxdf0bgpVrsoAU/Y2xxds+u98hu88MJ0n6rXgdPoMDGLt/asHz
plefSd0zeZv5N5nNIymLNDEEMoPpGpIY/oTe5OPLrPej3T6iEyFovoI/TyrOL+HgADaxzDwNgAe6
3CFWeEdpyRNbZRkGMsSoIIdrJFfsmKl06ZvR41L5M4aVHkbRVzYty21oOY9mAsYT33XzV842HLtr
KOzUHgkehtZiKYIb9bTxX4cmNJOLJsXKqBcD5sgKM8lo7KJEsqxLMkZ2RVyUx5HShRdjPwibi5A5
+Nn1w02j/Up1FLXg51Mr6BsCTUbyDR9UTfKodabNbdTd20NqbDEeFqBL1EuH43FZdA30IJ077MLW
uGksBVLM1LRvG8zHx3epo4OXDh/EseFkh/qOW5teMCcOZGc8i5hzFjXqZN2jPiCNhOinqsEclL/c
Tn3QZHCrCcJtDCSSmGbj0WQ34nxAA7CG2167jemLtapRpENT7mcB8DyMCYyYpIYS+bp8oPaWaFe6
NzNnAtnbsuGql6qXlmNbk3/+1XFTCvrId8v+qehfm1JuGx0+soW5BaWxvJ30g1QNhqae4861bX59
DX4pvzcTgIzatf1cYmuU0ndGolGLDgGwc6frlNvFw9TfuWZB5Fmh+JeJOKhg7H4amthZIBL6DuGF
kNh1NkyBOfKfHULnvlhtQrDLQw//VCnS+rX5zAByglW9aopIycQKwM6kLun6QxRv9R1XbC5EBOpZ
jrSDxXCzAXLQmdEPLcJZR6lO7mfqWQWCX/rpihU8W57BdXQj96A3hzzlZhZDKVtpJLd6YMTwocV7
az+PRLzQRpH8rZDAwQWHadeVWsBSJ74FpmDMHt0vzsXEfbaOhr0oIcNe90MOEs9RhIKRXh0WXyBd
tfkZY8cCSZu/bWJxtEQFtUQ+u0SuKSM6dmovdaef7cE8NBxglWw5uXXMz8EGV2g+PLVK1vsXnfp6
6zG3b6fHQFNFY28J/TeY8rrh2KZhD6/+LsIe/3WTkM6seNw7WO0r+xTBaQmmnATnH5qvhpBlg3Lu
THBLd5mBXGZ11FVPZuiHCh4qRjF8ZJmxHzUJyDXQ4q6/Tx+U7oXLlxFBxyKxZMpwyFIrlGbSwoBq
rZWTGSKUwzSisfBneWh7vpWYUmr3km5sBdXASy4zkqIfMQ6fU/obG02kPMTAFzXhxTPgYOK6h6sl
FEnPjk5fq0oMfIP2tIqKCSuDqfdLv5YRAMAUcOHFyA3EQWDzaGZzLLpt4nH23g7qANMDgNWoDqMD
qzCMcMJUDpEFv3ojNGDhv58qVqaDdtewhjwWf7brx6d+z2yqPXTGTE5HYcqnCWlmaXP8XxfD90bb
fwuj4CAEqzNSjDbkMwlk/nfa402R79tNdikNANENX16951F0Qr1xyMv+oZkOmJHYY6VzR6lzp8Yx
p3K7AEMiBLLvjxUZkh6f+WS0lUhKdbxQkOEt1xMYOHe401L3LQ6G8SGeCy+xVdr6Wo/T+rmN8d3I
d0xJELRDftft5sLvGEMlRFsSyTUMZZPeixKmJp8DDe/xDhCqKofMkFNJS/BG/ixlknjJMoft+HUc
jSZH/qzuQPJtkeG+ci8Cm+kO8achbNz/Z2Li8+FS8IIYbJkBTHP2/ryoRbe5LFD9rqzoHHHBzb/e
XzVUPZ5Hee8qLleVwK0HdrLIjv0UUrX7sHEnAysaP4mC7QT1gG/USK+PLyTcQjNJFcKlIjHkjMoh
iiXLXZqlbEvM56Cfpero0OEBAo6KURKF3/ZykYY8Ty8j6250eN8s1pRY+EzlQl5A5YNzZ+g+YCWD
kKDuRhQ7tbboglflb8KeyRfUfasLbqEzwyUdQEZkaeTpphNBwGGn7Da7OnWdmu0ewaF7Ys++uhGY
5LrTz3y/lsU2ZffjmYBR8ja2W/JIxRCAXWTslw1rs/jXkIRLDlKoAZsve+uCumGxLDxSkFVKQhuX
hxbVUcoVA3mNpm7Wm8qUfPxhiED/bMwL/s12U+9r/TmRCZelUssh6d1yKtGF4clUqH3RN9DboX01
m51Hp7TOkTLV1n6awqW6Y7HsyB6MAB94VVSBGh8lVQeju3bqBnOkbie2i2IM2jjlJHhWdL4v6kT0
r4Xp+2otGupbsRxnw0lp5GgZr0MqnU+bmyn1NJIhBCFyNakfHBEWwcwhtTMGCDQa/PKH9p2AyiQu
ITI8pHRPFgiPsxxuBQXvGLcFGaF/Cm8RHoFyVUVjRx4BhsaPxOccLWjdkMC3MysaZn5nQoeIlGcR
ExEZbB/5GKrlB5Fuk/PQWsaixqW+nRA8deOnaHdUrCisxpjHCL+Lkr98X+8bdmcI1sfJE1DMSiPc
V+f5yhJ+WUravSkvDv3vPoz7Qj1wCVqlAdAyGF6vlGIm8tpbdZlTl7o+myfU4GvGrNSJ8GYajCeB
fE78hFZlOB/vLLtkt0oYjZ2Xzd1mTXi1q2RXIyPUZdu1p6MODBnchuwObA60j6cvP+uS1SaPO+zO
ku4qHz9X7LVyIgVKDm+OmveGwhAE/UiiKJHR/tCNj662Tsl7kNxBt4G091Wd2iV34O8BOwecFSDz
cdxknDPgpk5P0KYKz+DwYiw9X0UQauOO6wUq9+4URK0HrssnsEe4osFGbFgS9taCbNcC4aBQyDQu
9i7C7Vy7pc8cirq9loWKcLxiru5DDCvM669faq5sBymQZI2H/bR9MmQRV6Feo8Bjx+DD2dS0ZyY0
C4Fw83VSLWHTIF86ENRtLQMNmk5+LatirMFtKt59PNw6PO3jQbAZQ7njLLWIrcYl0Ay9xxFVqo+I
Tbt59mIMGrGT/WsOMG3obh47+496pSvN3b8z9GDe5N4n60xD5LGJyXvzpr0DrEa70hFw3b5ZIj4I
c/Odq3d+e2veN/Gl+lrdVj0JsFI8PJShjjmXzZUpV0lv+sX0Og1Dd4WEVPoFYDebD0QD5ZElYPSE
fm8mkCRs4BajJoaepSx45V97LQaWKWJqYvGewQX8IMaeFN1hCWfe/C2Z9TjscJtvSfbZNQbtGj5B
R97GwLJrrInIJDLCOJwCsvyFqt3lemR8MY0n0JwxP5178to6KCINrAB0+mDztGaeyPM0CsYWRzKO
sxuGV65VmKySNk6Sd4vgXB+4jT49SxfLizrxDu1iXq1HUkAVlYjvruEmvQHi/E14Bok08IzMfKEI
y6BesKNG4got3eTHrdbybeqJBPzFKTU4J2DhlfACZ3Zqyy//O0PxRIZsjcd6c4ZIVdgBAU/hPawb
btEpXKl/MqDSPMpjw2RVpS3+BvTkmu/AxSNz0arZwD+9R25DhRlZnZZ6iKHWz4acoNyd2EFsZJS6
40qJQLYwF0emHOPKbABdgeOeUZDZZkjkyEDgHcJO7oV6txtxIwXvvlrfthL3g2IqO6DZZUaNsHCx
DeYcSWtJHrcIZ5l8HimfsTSaH+VV3tSTU+lEv8MCkiGov2ARciGkonemLurypRwAFrYILbdJmYG0
r8Rvi5fHueKAJNJ2Lyc//i7GOluMP1qRfSeoQEWz9kKsx3J9LQk4H/2SC2XdzCWjpbqI6wpPNfpf
haF39oIuVESAV3HckfMfdgj9yfwArh1Kq+mBGkq25rlTGL32d5M8IdqiZu+ShifZgPUvHNTiXq/M
MEZpyX9mapBtU/Rh8WLsryULV++vCcmqR271309CyCg6YFMYkNIXRLsdxEmIgIdTppfg5M081qsj
74SvAK3+FvE1G3ZKj4317QTS106o2utd7g3mKFuHAEU2+SDDmemOHdRgVuYWueTqBvumiXEM4TQa
ToI8NFi78olhDttbpLxyUeSUbYyl9Aq8PjNgGXRIYDreQMgg3WxjmPdZzTzqbd0WGWIkTLfIQ6GB
poVceKqgaHmI1WiO+7JXGEFzi63Pw025XGShHONSQ2xrOcXWrSrebrJWVxIUywAgpgbwhxhnJoUP
rGAgF83VK6C0H15KmZ0ZACTF61h7gepVBllcYbBNc9scalja8lIRVWIezGKdwMPprCpvp1hQ9jjq
gYurC9TIo5GkoXJX2IHCWsLRqznoJu+9z+0IpnMjZ3v12T7qV6GUI5tL9kPYDIwDF6y9gh4ZG9Cw
a2h5esMFbyFZdDSjhycjRMJjJv01pqogeT1WsKQ27QT+PtseJUM1ZnQv+HbCM0Pr0EeXE480++Kn
5GVYt90PspwTAzJwN+ezNN7z6NgIauNM1xA7aewboMoee5lQ6VxPLJxCj2copVXf68OCPW1isYH3
cAESreoLuuvlNqRkKxNlzwlF8OyNzkwjBLe+y341qHRtx4y25QPmMc9O7069ilkkdWmnqzgIa39x
Ztho1wJCc/6zRFGJvXgjdhFAi1MS4JOlRe9AEuY/vUgvqyBRQuJ/0Y9tg/poF0nhW4ivRca/qrnD
JRRrxZ5KXuyxOuROjBN38QTGCt3pPxGHwXmq02HoN3+W5vKGIpAi1ctZ9nM2iZ/f2y6V0/AzpPVa
Aetw0jObvKmVNW6wnMUib2HLQ6QsmFuK419Nw6wUMQaHaMncXR9c2EWQwqdCgfb1XjIZdb+SstUY
FoKRFndSE5v8Tx2WeLEreeSsJT2U845DhcZjqN/qZQOnV3nsPpMtm9pRxNKAR9Crs3VUkSjq8iM7
yzfX88XgeJEWu/FK9DT632NlUZbozirwiNxn2e8+LDB6XloElmnTP4LQ5ynN3VOIHbw3rtmi6JiK
Ja7Et/kg/57/5mWRgyHA9sSFDmXWwmTxLB3U2h0Ps1tX9XDrgq/AjYXPgXtERN0CmjBCc/gVApgB
7wRWXLREFS4hPyabAWAyR/njbo4tZ0wWzRM4pDOMq89KF8Y8rxMsE3SpNNPF4uhWeO5XxmzSQJFW
INEQK2hvJMYKHWY9icpU8uGrnSkQuykar/6y942avQeKANuMSgkYQa1AlB2B785js5yoi4F8yEnG
uIqBNHAwIqG1uHq46iEkFmnAZQBR6Dl9ZFpfE7NF/mBvOx2GlKhKaAkt7qGU+61iXHDm70xYWYXI
FNf1FC2Xy+7AuQHKmwkAQEwUe2ZSldfnDMBRkNrFxpYnLJv2BBU63zqjCUbBRMky7CAc8hpRCcuE
lX85iwWQGDqAxXGRCO8IyAQ0iXnL5EXfCh5Bq+3Z5e7JSDhvrWnR01uuZds7dFZWDe9B6Ld+j7j0
qkEu0HWmsKdlNkxBmUfXFJ8wFT/Y4hlaHlYgyAjmEAbKxOEcaTiR+qVF9Q2hdYbZsKRJMpLgNysz
XCP6yPrGRH8wgZSVX1LFbA0f3IbNtKFL7A47retXyUEV7s5+WIlYq2DP3q+4Xsl+CqFyuBkEAIeH
4uwWpPp8akaUBf+uIMpQO1uyRY0Ndenj5rMqA6BwvnZcszDweTBQ3OEnn5qXIt6qdSQ6mNjCenLa
l0aRsJdRsryWPQxoKd9nDBK9rcu37+2M/LGmZRrEnvo1B5UYqavjWwI9bY8MVaEAaAYSj8ae3cH7
nj5vIvOtQH0aF2ddQefVIbHRajHxaidZWYJsn5o/3YggZDQfiwRg46nh892Ism6iW4VJusPMAJk9
SuD0tBDKvYSYhbYkfOKiEcwJsPi+0rHFq7qVFhLQ4ti486fNcR5hSqLpYb8SsuxkhTimN+17ejCB
eUcvebw1ACYUxZItd8cNTd3GwKN5Z+q60PpQ+lAlqVOKkxzUXiuiLOeQalS4A4XQaDRYqmBcRi4F
tdDZK/LBPIcuh8Llq5qVr9BSEiKuGnuaWVtkAYplYW46IbZdIlAlK4J0MwN+kBakgkafZ3CD2ZQh
hS5CeiXuX0c+cfAQ1uDKkcUBosE3gUZuknRbG+H5h9Fq5hqAtapuQm/gQ2fDhuecDzWTeBC9mQj5
9kL/RMj7F8T8Cra2LhYBgLYmSFyUtiZoUfkRFV7qWEDCCie2Jv+YHEPECiNNsCr3UzjwDpquyBsL
Awcf+8NkvLuYCOlwDV2WdyE+b9as0jn5ZWt1FBocEsTGI7fq3oKt2mx3EXGqV0YyZHTMIw3c1pJ5
EPySwZcKgd1rtUDtWyX2/n1EpUtKaoChrtotxkr9n/YsDsmSEJp3Pr2I7g0oTo1nmkFxHIRVK+p5
3/5rVaJMRJ2p2M37UOShLgjmu8mi86z+ffxWpfAWRXCSma17RiWqiWHthrWn+1s5RKkl+ryE7Gvi
y01JqBMCztkm6Lw5Si5qGyTNulJb+UIOuV0xG5QC7LiuLkfYLJxNL8UnNxKY6kxQUG3VqaL8HX9n
ktL+70TF8O2jNsiad9+jDDWltRCCFT/V2xX0BbrCD/GlCQ9lWtuItpigi65A3sEKaDpUlrvG4GOz
f3SfDcqgpokljKw/gew4oGKQl/Rj61s64/sSKTdgAD4IA+HWammmWmmbbhNk1HljQGTv8JaNneR5
G0f2CVRKuGH55JsnVTJSJee25PacYrke91GUcZS92SxcLBDmo0Kaa85PBGKf96M2ncBXzTAsF/T7
VsungC/w/aENULYrdstN306ANjg2aQMkd2pluxYxsNBMmxYr+imWEIuEEbiRjjf63fMOOuHiGbd7
hoPuJLJqvRqwpR1rEUT0n9bVZvnO8KhkRRthlsjEV3nT4jyxcCV521GFqsaepqx3nj5W0ysudqyv
67mNtvOTeRMo5qBGCufGGmh+PIexdZv/M2l7CxFdKgO8BInr7FoUg4WG32KGJuown79h9bSJeaVU
yFXObpXatj7EFU+Nge0mkbKmnR12Mo3EgEwhEz+sOXNleyKTYBcY9yUiAIUKoCLlRsDxul3CJj3R
w6hQ9ryZTjH5COiaTbHBnLvcOqWOYyY5NudW0Fv+VGeEeVMrxDd8S1MNgTm7skrz/9fG1MX+9UuQ
nD2kK8/0ZvFnmCRlLIQv4Ibf06oSbrU4Tnm7FDPGVYjFh4MqZxgezl6FBXmja8Q1qdPCiduxwhee
3xxjyCdBbFSE2uLeoAtCrK7ih8HgTlOaoeZmXawcyjO2KdNBMPL3B1mohOE7a+wtTiwBhaK5/WSS
uZhgRf9e83PZw5Ank+FJurUmwDgQG5gXRwYhr1183GxUV92DKa1JiImJQAIaEK0Yi9o7YVHFqPd/
Y6relQnwRAEAnqAaAHzk3nntX7KXPFmdIrkhOw9ICCh5qdVmu8KP/y/devz/G+EpYMp0nsB3uHSh
RgTHyWNSlq+vOJo0iC2SVgE2b5moxx5E0gXdSixBHNG4TzPwGfgiJIDcMAcb5J6FRBhk78N02IVB
8IVTLj1D/+kyt3klzXrSavUZXl2ZuWFg0AQu0exp/bduDPHjBXBVNurm7xB14VNKL32SjRF5fTAH
PdG6r20mJnBZ4yEAdevyMj4Cws/W+Sa/K+ofkl40dOSZJ2ECQDlDMvZqj6dM3CHBsjDskNEWW/VW
RA30OOSMP6bSa27qeT+RTjUXVE2ATrHBHFTvS0CX42eR+uPmZ74u/wy4R0uR3+0+6RLvkcXZ+WYJ
XNKcGh80QVeiEhLh6Y0xPnpb9oSjH2PJLjtn+1bDxUiav+uN7GucYf8M3vydCxI9iuDzrPhIj1SQ
VocZdYdeOfIAYYj+k2U5BBqeiqi0Ew78IXMdY+U10nq1kdTTP+TD6rFarNdiuG/QQaQ1OdspF0Z+
EE0LmiC2K/gDmsytQZ1JXhEum2rAo4ReUwsowuqWTb53dzxcKzr574kxmpuWR1drL1GERKdocpfi
ns05GMEzGZtm/SNLgz2a+l4St/wkIhmNwdSOE6rqlh8vdybxsGbDMx4Fo0lhSGxn9Wkgglxkeq9c
WIsNFtR16R9eeKxIV7WPDGJuRb/JON3MEFSoq+B6iLNXPfOSYILd9/r3WPkqLJatu88Eg8CBJsq2
taXIxh/6YIHC69k14OC8ujaOEKe0T5O6BNIFodwveW7eoVfROR8wn7jF0R0sgdD6mOpUuJdesMDc
tpvZB42DulSGm0BGgeQHxYWSZ2cXIAeC05c4xLwncI9qdgY0i5NdVxrStqNPK4IB6W13G42cxkNN
j0KV9olyOEL9TKK1ISIw9lC3ifNGoQ5fVDPchKBmfjP2q5yO6ie0O0rgY/pY+aVPUIa3U4q8uc1g
PSS7m+6dr5ptcPlqa57Hb8tOVm9GsWmx07cnmhwRB12PAOkMWwN0MEh/QtA3UvI5Aho6vTRaWUKr
R9gz9qlVXkMG5XA04QZPo6i5lKA9/7GLD/iWypjgPAc7AsphfqopAMyxrQcObjRW/r85hcDMkKo4
lIhx9zYDPzBqNnyKSYLtD7bzoFovNHorM4VKKeEeVq0MAAA54oNag90DJkuq03DmdiTg9HnCSa0h
/PLOX/aAi2ZqGy/7ParT5I0lc5DehchSegneaCnjVNcD13X9c8dbfqysa8iaQLHY7yC9KJPCghVr
FLl/JJoGXxNFtvFK+UwxkfxyY780zN02XS/1w6XIvDXh/BxhZCwFRGES5HAvTjYCe+XdUJkoxTI0
TBf71Ze54rIGSOjRcr/wjYm/ery/yM2rFBKYQ9+3ZuPoJNmdnbtePBU623ZXUYu0cajCg9p/CEGS
OjscpeiKpLNgSt1S0WFYarmBid4c/EE6E1ol+Eb/sMN4x+UqOFkKgWc4j4ErJ6z0tdjy31QSBSLS
dflX7SrkKg63enU62pz/ECoRIZ+wayrYVs+MJntP6CnMlmLVDol5VHhRQBrDvwnldLUCypU0pDoG
MTSM9dgzzfXhfb5aVxNFu7DIbnbrsKFiY7P5Ru5srjDx/cGzstGPPaqkB2BVqXftPam0RoR69nR5
zCXZzWa+VM22M+p9nTo1N4q1I1aQZs90h/HlPvI+OTtcJJojIhR4TZaCxVPo2lLcxOQs/ndXLk0+
bFYrL0EzOlZGOuvOJY9DpTjySMuQPYQkwjVgqrAAU0nA2fvdFcYefT9okdoU6P0Es5Rl95OhuzTm
0DQo860uWFoLi7BkLDLVXHWm5LxEg3PSs7wZ94TMghMEurTPvFByfC3dFQ21c6jUaUbALev3j4Hm
GEkyOjBZYbAtMTwP8SqTyhi6ZObLd/cG2bNHLKkP++xV7xCH1C4oAJodIlBMZUJsa1lJeT9MCmhJ
qnwihWvPUROQIwsZ/Cgd0bbfQl2IUDfZ1y3hwQSnokowDljb6OZiqIMCWbOKpthy0OWItpKBluvX
6GVH+XdZ7UKmd0wQcfcYLarTuaUuWSpfoPJ6mKoL4RAhRAklMQPsu7buxD9fbJCVOxc/961AgzmV
fW67EP8rUfpskvNSfERdTFHe8iZKc3ANzzcTgTRqnJATr23UZ2XZzYHkBziXi8sPKNCPD+5YxRV9
uHrDekLh1nl5H6v4CZgpv9lb1HyWkaW8/Sc1b8fwcb1tD8ywAU9hp2pSc8vXed4k7k55UZQ5KWb3
v2nIGntafyW9v20Dvh7KeWVoSC6NO8gKakOkANkXt+pVbKAnv0mF7aLky6iKzM/TLNDnUJ3Nmlmf
PrY8HiBZEsAkNDPzD3cjGcs2Y8ZZ63oFuLizZL6cNhlvRPzXiz61RRFL0H/IjpidIxDnvztTlM5n
I1H2BXPLSjPxWYjz6LoFFvNIWBVV6jXFlHiJG0yoiai6Hz6tVVoE03QJ15zuV49tg2wIw50XPYK4
ckZAGc47S4NMe94nBpdxs/ui4XWQZJtsz6tUYztz5Ql9DltC9B0yUqeWyL+dUaUnflWNxwMdlEaO
07+Hc/Caiez+WCDwxJDSXu2R7oO1UCD3MOnKYu1gqni5yxubxQFJrT5j9fl7k8HjOz8dIJdZ/ZK+
lsszyR1kVBDOZTpxlPGs0t2HA0hex64MfbtlAiTRNQ1un3jO097AGQh5aS3/fGtgdZREJxpRPuaa
h4vmLflbY3oqPNbJWVCNtednuwo4R1E04wUwhfLVHoww7u/81xpl0tPAfnmwTDS4PaFrBiH3dzjS
YcQsQAlJ7uJNmXwpdb+Wh6WBeEoEh4IlzTWXosufgSJDtWw7jF2rrbZPsa447fEWLWMt0aBXAXNV
JhQLiYsDBd3cdkAYImd1csMCcOKx+WxNH6wKN3Q75yOmyRL/HViC3Bfh3Rlq3nH+pqc6m0lndmDl
CF8TQbuOW3lZZd+d6N9MFQP+kNsgU5xginsdeGDSC8Nk8ub6HY18wpPOwtPxyljHYoFIdxH61nXu
18CjNFc1Z8h5y0ZenD7frMv7hCiz4LPZaR42eICScNUcQCfddxGqTVYjXFjNEdVPVF5QnkKzVPkW
N+ORZ7zWZPROiN1TMCnt9+l6WuVmzDVqJKi9E3ejjMqhfHrfWLgNs8F0MG+IXyS3B43889pcJScb
33CjaYCxzeR/vAL6296pXljCTMeueWQtjqwtc+6LouLDGaG+Y3StnhYyrphy2zQj4dcwF7HVylIc
Z/kru7U/dX1XEZBBoz8lgG0scxctCdMZbBsBYqXjZn9yg8/ArgX+sazhkKjXIJ8di9MPp35nT1pX
1eqgbDWy4a9970zMxIiVe6b9wDIDwcIeXp0WBuVa6sDRLnfLYLujrhqFI5eXMj8vSf3m0gTwSCLV
h5QF2zShm0g0H9Qv6q+1/fXf+rU7FPXe5KomD32Bi5h5jQAgFGx+tHogp7xQ+SjQg1NZfvZQmESM
1jZ9F56C33hOyuAKPkKPHojWVj/r9JTJLgzxyHouyPBYH7v8EoqY0X0qPhcJPMViHKaMLBwG/yVy
PSnoafZ+k39ldMAclpZKPzJjRXMhCg0QG5mz9V0J1hly6hsl2pHOX5I9u6yN+fKQ68b6ribuN4Sr
5LywjEfEAKR7zq2QUsp/UffgEw3hl/I15jug+roNKX84h6Bm+xJ2VCOFhsnq47FPvkuoaRN/2vSt
6C0tH8p5Fn+fJqXgi6ZGr31+aERUGCkVsmM1DfrhAcMImMD49Di3AHMqjOMAcoyQAbplXPaPkT4G
ROSxD7C9CIpApq/5jVSDnkS5uCWDfRCrlW0pK+gf/churFT8hkxm9Mbu/yx+g9OsKUN/lX+wBowG
1wre+3beNWnxyQDW3igRNZkubor5ob78nj/R671D22UDqxm8bAaFpONlryPPi6WsXAVZy9ag0AtI
XxoghHQ2DGbBO1+OCIcPwN3tdqfxyu0J3uthCSzEzWyrbJcBncunmIRmJJEfUKD/Zixjm7vXa2Ra
BWY/khcOaHQDYjrZ0L/PTAyFzMKTCDMeBnpNmB1SbHU/8cZAHHPcJQNLxENx6DDPmVLMs5ud8ACm
5gWuHfWkVyH+/e58alq6E1sCPL2uPzHbTnN6mdV/uJj8uEvFhthgdkhvfvIqlDVDkzRywrabhOYH
dEwN6iLQSPds5UGGgJlXDYK1gcvqSgyzwV1xq1gTMML5hZcmFO6ynhsSP7Si/7adwmjxsWs0Hu7K
nAftFKJ52IIAoAU4/NACMzYfX1t4DFcX0D4T38Rnog+hWeu+hEYXLk/BZj766dyhr9gzWjaiMofu
e8kz98itCrdcUftotrmfeEHu/lZqevMbJX6TlvbvBHuMGjWXA5Rf4TVgdyzFy6K+nk2yaw51v60w
clqV36kDOW6QmAp+30T3ooPKJjMS5MFCnbYKrQukVRDaJHLGwEXob7p8jCtrXWeLIK5YKbxbUPdR
tqOSlO5BrudqR5kV9Jv1RXAexJlRhWu2CpkBh2uwrEIFynihNFpr25q8ekyZvY5AW/cU7OU73r1a
upSsWhlM8PoF8IRdslzPFktlwjvEh7+34uIDWK4d56242JG5/02WQlMh+ckKw+5g8YGOA1TiZXsi
tyisDRZgs7GNT4oHEW98qk0QPbOWIqCcV7YlqpuVYf4AJmCyIyVThc+n6upwIUpWgvKMW1g+K5MW
UsVAK/KYtDHUPYWS/jxZecn+7mwYxRTsFlMJqm1EblUqcz+wisVPp2GaWN3+mgfcnsek0VA8lU95
CmKtdSnOGD370oW8iuErQJLeig1BHWMT2qC/GWCWVKx7IMO6RZ69tNVCw2laiTF+LJbh2gW89kSY
UGLqu2CxABREwc8Bv83WBND3kf3vKoudNFypDnhQK/7jGkykII/GAIPS27jsH2JIvHSc5l1dcBe4
vfYFdrJ/0a7PpuSBOxvfOqSh3olPCud72xByzDUi3yQNv7ApzOOvKzOepcTANFgFzaIFoy0jZLh5
MjQRCrmpc6VQpeJfHY6t3pb8E7T00N5nHle9Hs5Oj6otMdifmSc0B+Dc1RIJjUZb/E5n7CnzoXry
1Qy3aeeJ9iwVpCBIzEnSycAzTwuRYRW0ZJKokGc+TuZrJrhMxti9UyZDuYRPuBez3fsvR12Mpug4
unMTa76nWBeCp5CP8MZ7eX8pHjiRthUfTwR+mq4I/C7m/pwlI2GeIwRr56EfBOPLVWyFPYetDWV7
FqpraHhTV0fA9QTyn+PQVGk2JZSpk7M5EekR5/1SbF8dZHPJW20131w7QDYYvMBcpqHnOKjxFova
OSKB2ILYbfszRkrqZcPNuxOtwZ631lumqajaq6RFBX8/bFWd6/UN9jaDqJy4fblvzOmccg5nlxxH
KXU+aVHZEKIy8Q7rQNu5FAyHF+U2hjbeDufwPrVwqOQMn6Y2PY7/vC3sFj25PnYsnujs0BGkFWi9
sdeosmbOQUyObg7qjy7O4R6bwnQkOG2zq/fG1lyrkhBH39eNk0JEWVb1F8i0HQnecJR6OzHcTA0m
140Ts91Ub/S3FiQ1wJhAgRpy70TH0x8TpGMi/HxcvnMD8R4VwlK5j5Cr8DhxQJ7la/4WTdLi2KvG
DE/GlxcQBzntFAG1kWWXW91C24G1whiRns6FtMpMb+WfJ0Kj97y1yoiz1x0wvSBDb/a/P+v/9+wj
RdDnzsVS8J4AdtygdP2/FwhfperbF7aqKdGlg6FD/iEb9awiWLSeR17kP5rbY0rmXyDCVwFzxrUY
tlP0RVnUKioZvSQoo2qpY7WyTmvTw9DJbOQ+phB1m8AyTmLj1uE7r3P2ZMGChmpbrym1SI2P1XjO
xosz1K6v4gVkL40yZBi2vq+wXQZFoG7+VlJ+GtSnz/rXJG1ysXjQc2qPsMGNZbcJZrkx6mXUPavj
jVeomkcIhXasFxjDPyQBKqabHBsMb2+K6u1/9ga2OHTYzw/QDIuPx+5m5/nMVPKRURVC1WdHwINA
+vhq1+xTKXIWDWu5vzZ/kwzR5sY4F17Wglg8Hmtr6XstYQ1Ph+O5zKJ0sibSfXgp50AvkdYWVHaQ
fomfFv/dQT5Dn4OR2n3OONdknESy457SmjysjQBFHhCxyscL46zfxQfg76Itt2ItYtBu9iWt//SM
lHO10S28PHT8mOkJScLdbVmi/VEf3mEW/pO4RWH6allONKTQFulq8fYfXCsh77xIyKuTW72NEhTt
pf0dn3VbKo0yQCBVCvVFMW4xPi63UdzUETDablMpBGzrbSDGs34hpQ7/gPPv+T1UDca0R7L73OmI
E1wmWyXZIbUSkIMLvonRtw/m0KGy5vjNB3lAn+Zc8i9WcKheit0hL4SCaU1GwIqaT9coVoimYoQ3
UAtgxHvtbU26ZIbEwYD2PZST5kLzbN8TrZF9NwXw8TIX9UHdtnUXEI9HhNYTe940g2P6D5F2hXyy
4dJr2ILxpVXGCWGHX2BEjrk3/hxwrfzphtS2UfYeoKdTgDk0WvZOtcmYDOTefzR1vD1IEmQBnQyr
cjXqYSUoICBApQXonZtQD1upR5Jkv10qL5LVOmIe/fZomuRX2BpH77rJcdesa2HoczPViOib7Y9f
SHJz7i9IMLwotZ4OhpdhvBNbb2JEwnttPM8asuy4NarQi6T63uZFHHH9WE8mP2HBtxAEq6lWCOi3
A9lRpTa+1kYphXzMtfuzvUJDVRVzU8NJZWHsNeKVRyeYmXEWLR9kYzXcV1OTgbn066DQDSudr1/g
ooPciWFeu8fl+CMzyIlLPbwLK0wzYfebzsJoxpn76zzrY7+YbAqhI0pU55gGr52bGfD99m7oMh76
rrtyuMKLWQDow7uqdbrkMi4hbSxWPlYvyDYJxKFrKH/25tnfAXmMYJ0X5MR0qesWqZD5qctZF5BC
PLAVFoZlWtP6t65GT+K/iyAhN8MzsX03PccIMDQi6fTvzaqhH8LiYPCfh3JGttpTz6jMvhGfsvKN
YXlkTvWHxAJtrDOTvWKLSB7xB0cYLWYSCPtyPtGap2SoKC0Dk4fnFI9KUmGL30ebjr1vzPUb92eI
rMADjrR0YHKj44WBCEYM7thZkaxSUHImsRMDuaK7HTf1grhAlE0qaTKUptImgl/kvFb1tIA3JsPL
BQCtYEtkVgj19+4Zmbxh+Wv44rYO0ID3Ldc1ZbRp9IOPrLulYoxkvH3o7PWzFsRYClQO5MZe9w3z
cilb1ohyCbfDwLXM1ea4bypwOFZPagy+rYlHKOJRaK1VzZzaYsomuv2kvFSzitJw3IdLxp+hdWjN
7Q4Lj7bwD133YikW7Nd4IFx8J2ujcd+RYzBdJniYGMZqXFyyhRiA+WANgf98tQYyjFLGLGGyiusY
6LVca6nwuWppHmeamEHwk0xU/eOso55fo3dhvb3nmJ1PuBpdS9Wk4CUGuc6nZ93nyPbhbEKOXYLR
XsrUkMv1Yrp5pGZI175VU/SIi5CTXZzNT8qhBCvqAKO65xhfZiokqqV8PTvb00ezwwxWho3QCjIT
Xjhf8AM2abOCDdx7UWT0h7Xu4LWhntKQfeE5k4JmRSQRPGrazWhC5FlC11GvSQJ5FVSkDpe37aki
afxKBn1+T6mjYi2aZ1JE8Z1hjQYG5TofWdoOrmoh9pU4J+MEuZ0/OneTTXr3ksq/FXdD9Cy02ZsH
PLV8dlZORxALvdfy5dpjrykwaUIRjtyVaXmxif8pR14dzewNdGTVTeELP0etuZcx/CsTzzRRb5rL
RS5PmDpNZ6rPy9A++tJxCOewiTCTA/ZZY9V5CThOVecU2hIM5mAgCl4jwGEJjmWQrqLPNgC1qbiH
+xdEcnKjomwilAcG+DHqrmLFhI+fJndzLgfzw1w/DRiN+KUDw7GpUf+w1NCiIsd9VO8eQIO7v16h
fjGH063OpazuP5JxjQ+0RCT0DuxeO+7Yb0jG9Prau9F8wpmJGxvVKJ481hp1QGYv4X/tOYbQg0sP
O/3fQpKnnOTLLcIu5w+WKfMZ/42H3ruFXELWkin8LaaYXBfHH6BCiws0fx/BBFmAD3Q2LLQ+brwR
8RNDxaFYN0XkoSgdz2axjS3dOLX2NPZj++w8OlcmdR0O6+fHiSLAr06JMJRSxZXEKrnU0xsMJSIp
/koCpsq90PqAsiUYtc9/TlgAxWllXoYZXQm7cqqDPvfla5KRcPS7aCDGjJtO+KFd6dz90SAf3mpW
a00BJTc866ZDET6sajwl69mnXFdmUg8RvhIV5BVE20sPxX7I3bipHCz90Wy20tg9jAap4k9XFzEW
db5aRQxiJ1nViBfLOIaqUURoQZeutIuiKVodI5+T+Z1tcQPy8Zu7l029fhPAY/7QMWvKIhEdh1Bf
XwVXVpWiHNbR/IGKXwdOKaZ5ymWSyPd1qw8f4OaVinCQzaktKyjromGMhsgLLLu7bA94TnOmsRHr
B/EmGD14fkc4uoVFkFoA9Q6CpB0vfYG3RvfoB3YoBWreUQHc8Zj8q5iypAzjjBIN6EAsoRd6Fgd+
zWYuNZCRwmZXm9qmFzlXc6SL5zhTpce642lRSUubiZi8j5m0bQf4axvasldHUkgivjjyww38f1h5
FinZWYz24zLExTeUfrMt3ppEgyLFG6OOysjxc1VvFW24sqApexwKvBFGKAs+R/ND8ag5DgtYn/6Z
fEyWtcB3SaquyfYKAFaP7+LHXrIbYoY30KayVxWkr8+LD5rQTlvZce8zBLTAyUcgtzC6ZhpjXlge
xr8KY5GFStdXpjIuSyntZomsohx4FuysmCHfJsoxpiYNMtV6mAubLs5BPt/f35R4ZkEn+AX45bIL
Oz1iaO+ZYaW8ibTd3sKZcVG986XO5oHsXT9ZbRm637gL9U8z+y/sGm5Kijsxxnh909Ht8K5enWNX
/42jPX73iNbyCXg/Z2U2JTk4NOXEJx7WVc4+uKv9xO08ugMoktokoldEck22aSQyp3/9yusfCRA/
RhpIqpM1kGYmDT5Xt5tVOHGacufrwW0CXXMXqypHFfQ8jePpzq/gM9SONA8ZS9i9KR5dGFD+lcNB
3/4/8lvf9QgdhLrI2aTccGsXEJqYP/WUhr2wuBrbdYD1IA9Bx8zWg9z24dth/YoaGVHLqzh+U3v9
f1OKz2bilynFwba96oj7OMtcbD2vUfbpcJaLsLPAcEnIlBpaSu3pRV5W0rARW3c6f1J7OjNxuQEu
wyGfBC2DY/nfU0iUg33vQqyTeN8Ar9YeNllKhq/sB5jQ67N/T2934MZQCHJ7r4X8XF+Z5Kaabagx
3Z/Efmc0pGFuic7j91ApmNLmbCXtFkjxAr+sZA8GuqM0Zh6V5Kht5v18tAlPT6h/TAruioKeKkHn
u02G/BhkenSjie126glUe1eWsF8Jzaxzh7jUs/TxSsWGm0UPFX5Oa9bD+7nESiCCmgLsUojVHSYP
mYvichpXGnWZNgEdrF6L+rVilfJFy0SR6vnaeIRctEW9PZK+sPhLjC7hSeF+vU0npuRyhc1jpm5y
oOLTxBAM8paqlMl27jkUyMExJgCWt/RMqn0ikswgy2qI9/0g3UcW4yXUIl1omps+moy7CLMY2Mlb
NuEaxNTSz92PSLoxcp3hQcf1d4O8L/ybAKS7L+hsBNPloy7jHSXtqScupl3eX5HjDyQmdr6L3kZc
3Yb4s4CA2W547q5jBYTAQoYpyWAGyKaXFvdEdZ0XXTK2ibVzZ134hPAoIckLFL3R029hdltFyexP
Nyc5jzglQyPVYChLoCrBDlgjhGlR5Y8qUeaVmHu7rzhtf1CNRYxHBg5tjA+MWRiBVyhiWDfEtrdV
GmLBhvysknp3x/NGCSAFvkFe3vk5MZirgh0+hTJTAvaqkASKoSZXEU4TF320pm+lXxcFpsQltKNA
V84ReQNdl83NVubA3N2NtAPyTuegSZWUhXzhOWgKvc+h49D21JJkUA/osdDYojKazMsjQhg6tNX6
mz31ARccVVRhvbwWpwfJud6VRv6jiazsSdnTiWd2/SksvC71eyp+o5NCZiOraAW8MkbxNahR5frq
LQ1CHT8oT17/6L//CkiavashVTNtx3aSQlofp/zhlVKp8D650gDjnH8csNnOffoPsbMyPVWw9SLD
cExhX5voMhNzadY+q8RDLgFCkObXPHksDQrJkHDqiF4oVfJQSF9rAiyaZ+MKR7Hv6tDL5DaD1V0Q
knKFNAbbDNvfc20VxCZ8L0Dhtz9N6lbpIBT1ClgrHz3nC5G6E/g3iz7+OMd5rdQQzObczKjQbjYY
3GG3tHe08PJcguce6DqeAxqmzMuEsUFDVJL2GI15ZT45SRTKdc6iq8HBjfAkSvjAyl3Pjib7Brfb
eVOOas3ta2RtJ6ov0ZxQ9vTQ/7JCDDDK/TBgoMOqKMNEi75jskmOiFt2yt/QVwk1Khs63s535c8l
rvBJF1MpOsTNTQU2h3En6vMMrkn6XHHzQ6bbXvzg5OyBW6/E6nDC/DTJrcejlErb8MySey5LC0uq
HNPwDbog3lzX57aJ0+xqvWRuFuRdfIO6SVpm+WWdUZv0YB8gdP9Z5aozaBGv9guPGLED8AOJm+0R
9osEt0KjWsudoIOPDgwVDjZs7g+Umtmz5xbHPCiiPCBu6d1yUVqeQRaBFxAsfPHOQG6PTEEBctiV
tz0xV+nPcZYHxccHZYTlKuK1UeGm+QNhzVdI+HvmOyGUknwde4n7flJGqxMNjjrreMB5QJJgbCGT
ZWeipOrNs9wevx/9hQGppnN+01wCK2ImNcJ7vxJDStsRjrziHIPXf6q9kMsV5w5HPNExbngz+Ib3
hVTUxDiDz+mnsHhtZYrOUwsQPfDgQNYRZtGnFgZnlMik2H98Sr/Wrwkz9Cfw1cdm7jLsZluinXXe
AtV6YxTxdfkjKGHl0d3aAkcZB9Eo3ocT4oIL6eKW111ShsihonyjMOzyjOe39tGgk/g+GPMTBbPb
oMZN7cMDjYDmkHjOsQC/t4HbWtiDLUAoQSjK3pOzc4/QYmJ+whmlXPS7A1Ls3C35hikNnAXMRF/8
I+u9HSguXIiatL5DiK4nj5LRbRClL0E65ffoFv0EUlEyfD1KIKf/BdvoBYyhroVRVJhw/oHVBsSh
Qti32V8lkI7e9RFdK5n6iaVO4XUGrDZMzSAr1aMV5i4R4auSIenU9HRwxlU6yg2+72riZdkPXKr6
smySxr3qI623ctqYs5XHA6A1EQa54P1co8oDgprnmBd3v91fvTbQuzaUzEPpWtM6mFhm/4j4HYlp
4fgHzkTV/g1FXMA20TQELus2QFg4y+gu7smbH0+6oHackolgctnMpd/SuDf2n+IgnRQI0Ls8QVzE
VYsF0c+a5ERUlPVds8int5U76Sqw1/FJuhmZmzDtfvJkOi9OHoACziFmAW1+loLd0Px+/RpuGHBW
c7tGyUxYqkrC3CQHRBtzPkyYVSPe60JLFCQqYTfDjtBs6VzE8IaZOouddnz3MQJMl2usHeELM/ml
FGfILnxEqAGrkp85FrOfi9LpUBjKTcQikXXX2BLBSqG6tc9uzGAFiLUh8hhGHKwaIxylE9GEBCJa
bGsX9q0gum6anmNdkDh/nLDkSRURbkLRiX1xZJzAh46ElFJZaHJcavRCfGHuAWmD+hnm2vQBn0wD
VjrMbfCFSWRh0lPNVRfdQubR1htq1fURJiigg/lIhnEwABvNNYOy5ACigv21gPg7XiApyo2Crn12
hsAVl1SFnYXxdnUjwbMihqJSGYTbQRD9JaScs5wbXfbdkn19rxHCjGwHj+wBI89+9zLgkh7VhW7M
VO3r4ffDHTf1INrLsINLmN6Y5WeKDr9NKAhTfLmugP/N+XqVQRSYcL1QXZHdwgYT2RsBgDowdhhF
ya88w7HwFf9c4FeRzB8btttvBlYQ6Y2c/5EppjhMGPwd7abHJbOyN/A00fh90EixwZ0hSn8bV9Uk
CieJnQHO4Gx0Sz6F7JE+/dvxm1aP9KctsK89CLZoN4fKN8Zp/eOJ+8kvbbu0kUfLfFQ7mHR1klnz
gjiO8si5lEX/3HZQGTf7XVkBmtXeGOT3NzfKVuwY0xG5qGHKjH93BX0odAWdMdp/IoQlGGxn3ORs
R0dx1KytyH9MO5cp0L+5nAkUh1WB+UwcGSexj5hHMzbDz7ovGgGmJSIiWrAs+x3gYee6VV5LYNHC
YyntyvRUzmujp8B2G0L4qkHRYRDs/fIAhAMv6d0jR9IdHfGMpluygiuuogNxFEUCR3N+771MSlij
3QprypxUu/HidmDmOtos/vFtpXsxpU5zFclPUtQJYAOX3hykIoRowVZ3rtd2bytDXGA2unJv7ilN
IOMfbyy0ivvJNUlDAOBEGKC2SpSSB7qGWxvE6f/2DoNwXbqpWysCPP5GG8OqJ/zQIuUqpD3/D8WB
ozKwO1fOooXi9AbUH1fUX0cvZkFHedVIjA96MFJ+gOHMlk3cCHMZXs4e+1YBh8Ldiu2/Iypa1sFJ
JF+NIbKLUvZ6LhmUKFAPnqjZGb9VeFNyUmFCjEPkZjPJej+INSxVzrVsPNFmq9V+xDVAoKhVNdx9
yRUaRvDF8A6O6WKIgyFJrEJC20vV5ctz6jdnzF3GKlLzCUZpwXYL4ghOHNedSJkJq+9UTVOUjvtS
1r+hgH9XYulyzCRJPyWudfHKnLSbGxu7J3g7spYhQo1QjF8ht/6h0I0zpJ67numxgJkuWgmsOUA7
NmWrcBnhDE3p5zKULhhbzMVGw4zg7ACnGtROOkY1hyetHmhzbzHqRP0sGm80XkQSoRT8mz743K7N
DVTKM/tGa1JF109P7fRGeE34w3nbQjfGp16S7rDf38ZhtxZOgPdoHmoi9oDPy05XZygQhPSm03UE
NPFRSywbM5KRpR+nfepD7fre5ZX0ZuOjsLlpgaT1uY9w7QzhFWtK/QleONoDRt6+x/KllxnZX2n3
179o9x3jh+n0Qej55LVzJqtUzilkD2cESTajx/kXknB2KUoEB+37yo6KPsT8++9+5PGsvKUlK/Kf
PqgPgrPpAQyX8wJYf2dPbdqbloIQoR8HjH3fF7G1v30j1XT8UMj0g/exQzOoodBQVdABPuCHCXaF
jLihq1djA7C5QJMCG5x+Nnnq0QuO48ciavxfInu2dfypY6faymgPznI5CZxWexudoRj1jcHH0D/6
ndqBqBihaMmkWIHNXZUHXjQH7U47IDqHWpTj954K1cuHUJ6VrwQzd9zSHzSNvTdXV/sI2G3RmLH4
ln6iAwYwNSCRExqA+fmlSnC4py1AOvWUhwSHk2aqDxtcOcyogA+HQU/Ve6cLeV0m/g56hhkzQN07
qy+h9PptdiI5vgqhR8QYc0yVJo6wD70h0hZZeTl3qtM0E1OH+FB9RYaJDPF5+a6oc0/oTj7Er59D
LLgi4qxI48fGxztZfwoHekRJqf0lbjDgLHa/2Ykgm8r0fBgTrpgm/nSQIgd5+IVEuFQsp2jhBUgi
H4Sbj8vr6PJMAEIDM4RRc+fvWsF7fyGYxsKhpx7KxQSF36bpdXELuK2nI8GqMII/1t2BeISPp5VP
wZo/viiX0L1yH4c/Rl+LEfqAbVwHbbo4hz5DdL8Qws6ocdGFUC1X6Q0t40GRGo/FqOJQf1qYn+me
J5lqLEpscSSoVurhCOn3gM+bj/Wvqwbae3yztek5E7Gm52lK1MgCiNNVgEGiu1gmQofuldzvLArF
HDnPVenM50HrrbBGFyVs45nYJvNTR4tItabNJ92XkWwygNB/V6NXJyn7Bzuxv6DbngXyvLF8hbYZ
BagDgBgrVi0SyW97banN0dSiMoRXdSEJbOouWICSg7bWfiFgXhi2B/4EcQdxYOXU53kt9dnhjWDU
jpRupPldRRPgDntQTUxEooKUKajH0rsktaacjuVS9vmVqGsymbmWSsAHnrTz5Rt48AqCrEu7K7LP
T8I3XC2wwmBRhvsu4pfffgqJDqus3OL1XkFADVOOWiuXHpvtSDAEGEPS7EBHK624o90kYg1L5RuS
vM509faswqCxMQtSuJ8BXYrdp/UzfTkGQBvXDdBmpVHPkQM7sz+3qEABNXIhMrLpgfZQJzbWhv3n
vm/ZSPlhqszjHfssoA343W2o4j5dC4dNXrsSZG9v66pvtOA4tna9hBYgFuDinr+LGkGswTpgFAm1
f0Ri5VnyKhS3B610o/DR4io5fzJGq4NP/FqahkWkfCBBZeMSJZS/ua3/YJgZIzk1xDSXxYkVfqZS
bvxLwCltvqKccXsG0q0Bobhxc7rdX+1xq/auFexdDPFpY4H9YwWuVBbDhKp1Shb/7mF6dHJZ2sQJ
uspn4JqEtgd6Z8/1RtliTdr/2cErsXHbRXajkK2ieDYO+n3ffqZAbigePrpFUpfG4v89agResyFv
3NUxpiSHB6W5ohMCcYhpdCgHspas0bo6CMDX9qxoXYEfZkpIPBscTATYYaAeGnVzsBV1f2j3p2AQ
Y9A7qxqMF6zorVrwDZWtklqCN6PJBetoc2l/Nv2Qmgi3Z+m2B42DJQpi5XZEzUOkDsVL5pxpZbYu
TQt3QJOphVCSP53NT+s9CiNXOhampILNRwdVFqLeQ5IzU0RE5alydMWw8PNabI1xHsbAhBOvCYqb
QAOp3u88FF7t25GamieFml4UxNdq2Lkoe5NzYlnHOXODJ/h+DMiHJinszoXh6fc+XJDyhOn775Tk
ZfEBrtXENuafqPfjCKb/tr0omZB8UNaXngiFK8mlTS0O6xz+F3y1I1zxJrdMc5w0fUJUYnpJ6v1f
LdSut24CSRA471QtDlQeVTFse8+qATgAr0cnK13LY2mrMhVgw4DPKg9Fn417gNcHhpaDP/tVdMl2
G6OE9Eo00OXZqskHGcGYkiGgU4xh+6fVnQu4gwbt28aQAKE3W5tgFkuPo/18TzP5QFtjdzwaojZB
zOAzOpFgwc4RfxQet0EUlTjfOpxMEfFUd7zwDJ8dkQzUPM4SsV7YPfoDtevolaucPKhvkLTQ07qu
eI/5vyQvh8CPWD9Oa19jjmsKL5WzTsLuA827IOL8F9TV3T8eF4SVZjuVGJcSERUplwWIv1mymay+
1mHpB0mX55bhLdhj6UaT7869yuubIgnXbnpWZA8XfAPgZmEtjOGB2w15dAlGxizmsRsbp66eYvEZ
DoUnCAvTCWPpuyVEG/povXHJSoDWpxhRXEWwmrZVwuqK0I1q3zvLhqQKR53hmr646i4GmMdsYNm/
KSRVsmoivjoEVZYcRVq3NxNBG+Ez5v+MMxFVIwVt2zdKXJ57ji/LahXhUj291CTwS86koGSy0IrK
A63+lnhEjyGtTzVVqSNYaAlSMGnzibv547vTWVWpx7Ka9A3wMXMg1A9ldRjA2oP/BivgSrV92AXG
DPDshScgphNNJzaEU7dxuyO57cXkhv7WWlcmEngMMGmCi0tyHpsFbGSZaIvu+yiOeBxbRvImgyog
VJwzw5UTxTVM6E6BK3q8eCsumOSC/F4YFaN9z9RotFnt8XzZCddY4EoIHlyl6VtM76SO0/63QTAE
lCHpgTE6n595S1AekZ4edhJxIcGXsoAtbLnyyGhh8fknB+NugHk7idRMK42J/kRNUvqzrvgXOqQl
V8XyMRfriwf91LPJaiSOBpOSrEVxRLCg+taRZnJzK6CHB74+NIw1p5F1TP0i6HteuDRUrBoMjRQV
67JZLL2qQbjjs7hu5/YCt69GoQd4Gk8BSCYF9BoHpKYKxZ4uM0IROUol3Vxdb4UKEgH/RLxyRayT
1KjJDgErSWSkoglMbfKh6BJEliVXwig4O5ouZ3VLuDo3QiBrAozgK+kkfNqYMoN3Isrmto6MQF/7
9GHQ/1O3nMqAcIGDRT9xL7fkZ+/j8i17+DaXnIsyS1yq5WWGCOoU9Zpfu296kCfe92LZJhy4tYW1
xFW1H4e3TlF4euNyRiVGH9oWp33+sj9RUmOncrmKyojO50xfGbiz02ZMTcQjQ5RaYVaFZMBuv5AH
Pyw4bnz35JajnU6JIDzSPlu+9aDq7z0q0mN/a6EW+ncH9Le4sjztZQl3Kc574Z4Mp2mXtHIN7tdn
Csg33a3j6GFEim3JDTF3krjksJmopvFn3ysX7rjdjqToVmuG1kHbHkqG5dGKn4IDrbFoZ/FF9gT1
loltQ4zKyWe2LPsOtKmd7dJjvjVPI/DQHzL+GpH3KeUWUFjU9acKVpEMnQJQevi0TR3Y218u8mEL
AOOJN7s4j3SfnWWJKM0xCoBm25FyhE3yOTdp3u4NnAwGNscUy//056EiL5o8zmByZzgLeJBaqY9z
zh/K6lyil707r8hGtaOwU0vqhQF1x0TtkUsp09s/KyhBCE3U5ytL33PQsbnAIS2arLnVrHUO4Q/2
wbMIwLGZEVZjDCgD1Vt/mvFhVhaTjvP3CTNhVtkIPxp/o4ZVnOewrrrXrJG45p5TD1RoF6e1LWCc
iEvrCTYf81hSnMYsh2xkxD+CwvJceZEybCaxzsF0KCya7LvsOMFDIlF7ya/TD1ixlzs58Pvd7yCZ
Gp+gEhzR4ds+iBVsPxbSciBR0AZFjwIYEUsnkBzSWUkn63tel/Ig2dvGxJmAYMVfIcMlXl7WBlId
BNAjZHVMPVGaSPKBFTNwIEHahefbGYZmWuCVIDcv3jysubSlvl3EikjXeNfwk3jBR6t20PurjN8F
ljgSCXh/NC5qWMlb+3pSKCZ9oJ0uo8vImDxlK3qZ2H40396sYtNxFQMCYw6JFn7yHUQwpZqK21X3
DV8h+RmIYIKLJTBW4jlmBlMjz8tYWrqu3gObV9SW0MgXKrJrogwKm6Ec5QrO+WsZ4ZeiSfaOLJPT
G2krvv9lM0BJUX0NCzhvynfI/4RmpOyl7hg+VmAMId09dVmP7Sia94bu4Sb/7JfbfS8qjl/Eoio9
Q5M0x9L0lzJziHxxGYHVzjopF4cNe/Er36NCKzaNnhxBHDIy3S2ZHtvyJXOiA9pbuYtx49Zrq/PF
oamu6fvdOXXcSRBQdq/cxIZu3MKn2N4f4ifXAq23ZX/UWq2ysjk/NW2j8fvofP6pY9FcsUYO7eHo
M1bEcUTlulo6LqBl89RNgNG1VPr9PelijYFCatt5AVd7NkAFQY4vvvl9jPGG6xDDXrU9v5939dRX
1sgZv+vWvk/WzZKpHGFYbZoMaHvEmGN77oNmOcWUjb807OjndDc1+ug2Ulj7Vc6+JernA91jER+w
0UjxYvtj11bdvcz1rxEZXqOvKIyAQmFBFlYEYJLm1oJ9MKqUVrv1WNp9G8XxUEn1UdQ5Zgq7PtqH
L5sZtDlWrXj1fk0ZcbV+2tjy+wXnSSYUR9/4x1N/EcBtU9zrwGkDpiaB7qMnxH81JVKupGyUzlCE
w83KalgIKl4p7vl4MHvAEqDi1vUEFZbCdjw/53NC0hWlBvJQocNPLo9TMjmd7phvjanGLRQ4lAJv
J0IZV6+I8AMmsdcFyBseuThhkw+d0O1gHt3eVlDij/iKJ5JrjL16CwvD6hrpjjC5omvgXmEJwMdY
/gLlRcgO80/sVyCKgTg9kqMsPbQ4B/aJhA5Ip4u1PvZfi/wj2KnBu95xdDG1OM9n5AsKAuI/gSQ2
xDff7RYnhG2ME6L465anNfABDjKtOnwg6w1NO6RleLrP2dbKWzvlGcCv3/S7LWMH6nrogPABfI1q
qt3SY1DTZ5I2v0HJpPQEbqn4g8dx9VEeHCbPK8Hg1C3bcIGDeYeytocvxshfLuhDW/YgNJTaO6sa
fD3WfvflINeUCWAM/175ttg2vXUsBi8a5z/9ph0d6sC4M1Th+rdVdEXYkPeeUx2HAxMIAwk0SuLu
mJVOet7iDgzjPtNvlVdYTWSu8006y4Xz4lZQscpPcMOja0sx2CSt+4YtAB3+aG+cTHdqNew/VghS
jAyPLSRywtkTZLxtGXt0TDcfMmEhCPIbt1WfmOqb9U3Aobn6F6jTOVisKeOQ4HNyQ2CZD5g8J0en
5vgACiPwSNkaxZUfVvdiOcEarR6AwQS5DDi76rU6zVlQU9uU0vIFITRym1miQF5q672Rinnd7vKI
XMC8BKt/QGDfTf3HkB4cRcszCrRb4v8ZTDPf0KjaTYPYAt2yIYYxkllUXsIpqkg8Gw8xYQP7Jfd6
RKa77wWyug2hEjGOVZLGtkJIRTlrOqXHDZZxZXpfi6Td+UCouIwq/AVBSun81s2FuMUVhK2B8gaf
dHD9DB5Wc8/CKNcf5pDa/zMWR9o8tRuUE2I4xphNjxELqckVp0LQyr4p4ztH6S2858yfsfnnMdnu
V+n2ADiJi+vJX5I85c/cVAwwbscp5Csv+/u0PYIyxmn6oIfyXzJKZhjMSWsHs5kpDlizooXlQCBU
7Wrff/aSZVh+uFiKbZUHGdAjeXQBQTEhP1NTlaZlZ7OQwq4qfxDYTFGzS8NhM9wugSyLmCIeygcZ
EJTnvVU8UgG80iZGofkKi8+2atRoSmiERY6OATxqbnA+trzXgF2+KRjwN/P/rDXbd+XD3bg28LU1
DVhxcZxsJYavJLl5DEU7zSVr0pQ5wmAAciBCp/weOHmZRsn54MpdGq9amfvhudVYLBXeQi09gmIl
CYVHeH0voeDDWdKAEPY5KGBuDCRFJfj1soWf3fIzwB8H3dIAs1M0r5x8XJzjkejZ16buBzhtwkkY
7W2qatT2+XwQ4VfugUuiitPHzSrw09IrglhjOw+rDQDmQMcrcKOlJbUla8gVw39Tk2xytukG0x8p
RHmKfDMIz74mscH/BrvWB3VeK9RKaXH9TFGKdeNpqzXmPcT1N5IunzRHLmuymKhq2XQScTfrzh9X
qXlAT2XhYk+WU+KBX3eN6sifciK6RXG83mGhxo3aDQQbtkWPd5j5SBpgCoZSXK5kXc/VupuYz6Ci
o29SS/vjgZOb5CXrKFMCAboLyj3ws7ksknjuPiFEXkIfuHRY0IrH5a+D2b8Z2Bs0Gejc8bjlxVnn
g40EMystFxKRAlIocK0eLVv3fM6G8gcuI7QdQD5t5h1YRuooOksgp+6uep9XaUgBCyaTRDDAt4Vv
599fjpJvmP5gC/d4mk9AIbj2n4FSf/2Bj3DFsqEslpw6xsWcY5U4wF7lFAsV0sAlY2uggDMAKMnN
foXmGlrzrcDD9v+ZeLKGamAArCJP2QqcNNy9+Fwg+DU9JYrx9/FAIr1Pmbs0f8AK+8c/+iYGzJjB
YVEg9bHUph+dCoPzFJnSyrzWVrLEYm3Fm4cdx4rLFwqZoaMrnntvcf69b1Z+htN+HnWi739Zu5kw
NByGtXfGxCTi1pF14xTmy/3P/sZPeyr/hUBc0QW85oTluJvZzD6wE2FNiYjpcl246TwpgApz90zM
9uqOS28Brv3cMQ3IYrNXKiRXgA1hUzjTk8ZFzTdEMqrhiAbIXORiL2yVjU6scOv18OeX2r9VQ5JA
tttF0oVmqWa+Bn3LoEhnkb1WFvi5IGbWbzR0J3FKo29NnBiIA0vFZdlarDuQkiCmhJyl/quztNxZ
LVmx0r3L7IJ8lYs4VnpsBTEByef3vzgHSvOx5BlDLBHgUNAGZoF+i6HyhD82SUkeImhCEBxO92/E
BR+NJvqGofIJk2RARCTp6nHH1NsrN7oeAZ5P1XxcN09xA9SrEVcGXtwj4uycjLn/17CKrH0Eknbk
ZLk05NEtgEFe6GgPfc9w5nrrD0Gx4ELdzBQLuv0FuIXDJmdtItkecv+r2eeYaUr/plfYldrA30J4
db/62mgWnwK3SSFWVuTg1jEHhM89BVJmGgpG5MBDU/NKu4oS24kRRFKqxBpeJ9tD9KUfgUCt32SW
XnF00zm+AhT9nMp5eq3Zf0rKBsfz/ZhH/2nb+D7XyIcM7o3UQRk1Sd75fH5Yz9CAlzqfp98C6c0D
vUBiWx4IFPm8kMkFMsmOocRXbgq6yICUmVq6mpYKvjRNzgTtRfzQ9quY7YGxFAq4ugNZ+19YLCoy
SsFPdvLVGYuhdTtZH2fQXFVCLicrx8vnxKWF7I3s9PhHxPaFVZaTaIbdJ9oJKY3vCgEXpIP/WyYo
gZtRsY+vOE5wjqBu1+iYQONqiQol2zl3oYKTsSIeNIb4QRgafDzY5lbKadEikBZo2F0WEcY/lcMU
8e9BiSaCuhg3taW9BFrjocvFYRAokosP3iiVkGCjw0niJoRO0gOK98P1oYY1Ji+dsmdrAUf7eQcH
J1QvmLEI5srVC+yh7n/GJpYxnSHb4z7wDZiqRjRfwTrJ8XWHynUkl9EZEbxyYojXMtAngWEdufM0
/xXucTIcN6j02JWIw0XX0sNK40mN0Vds1KJFhzGjWymFcSEaKtNkm8bxXdu7FACQOThK5eRw5D1O
c3zzoo3MYCMjOnH+Zb4MYY7v1qGWqLiaYrLpOJ+wXHN5muDG5NddqQgOVcU2GuQwVpqKucx/alPJ
9h9m5z6Pz+awiNjwiLLaKgv3WR1PYy9/ZmrcQEzHCCzKLhPOzXvbcuGdyTDnP0UeVLjt8rOHkIXh
Qrjg+9izC2km4K73vjiKUoe+Pw3TYKgLK0JiIaUOiHbikHM8gHnCyGIJ8Dq+R4Cz2LLCTRPj3Rzq
PTZnZkgsKn+jx45GAIOHCwwFMfMEDWqYLZnxsZyNlEIGeubTsQSpUv5VCotPjFE2vNyxTMPkVnM3
sISNNppat64aicGnBWBPNji2CcX72aghfJdg7qmOSr122uHt8fjt8foCFARtKvocRVYUqRCPK0BJ
s14Y5SDlu83WEJ3Hwc9EPPUhi5XylcMicEIJ2zWyXFVvAYJWjMM2cFxo/9qAEOSgR8wTDqKA7J1q
S1a3TB7ULrmSZgWw81FNxKEN5GfykiD0XzgfYs/zLjBabVXoN++wbwk4GPilZNfASiftRqSZJA/6
Jh4mISLoKEnsbKy9CXWKiJzG5lNgjjkYUAGYA38CfpXTCtelyDpPviBxfv6cUCu2tEDJf6nQIpim
qFAsRm7Adv6oG2OKbVLC4+zZF24MdKQeFUXO/YBb1qzLivHYIF0NBzYs5sXOgMSPbRu4chAStOWi
EqnV0EqVq0J4hgkLD2YoJntksV20Oe2Gem6V65g7TQECSJe/fmGqtt5rG/TCTsgsNq9deXaB6Ke7
pkGLQvBlRX5SCnP7N14Z2QGU+ddz3GG1+I/i2GNUWefVEaxTuH30Af1Bhtxrz7qxUwQi9vuuMMZF
dJFUivVnSIdfgWUgmCy4ITr+cpLdJVxxsu352iABQEz51fBA4hC/pj63Psq90V3jnXqHnqJ5IbO8
CmNeKQV7mMSQ9t3bxIyYKc8HBt0GUAPJBhgrLtaMSrLXiHrZmGQk1PfXRTm1Z3j68wyD5WJXHED/
1kcWbLxfsbcXMEapEdBE9wvc8or066aFg7tDqfqxDdmZRlnKYY2QqzyXIt14xdsCB/PR/9VVFfIM
eoKcT+/uizp8EMMQkqZY5FyXI0CZZLojyvaa1kx4fc2jvcEzB2qPg5GvvWXUW7y2gNV2ZSiKUw2P
Ifcb1JTS5OTNrxhpr4XHwbzX5cK6arqzIBWM9eupSl0ats7qk7V3NbPMj+7X6zuSc5I44o3AS83L
EV+a5f775/lEbnNeFSPorap8wHCCozhTW2PdEX8xV0a1I1+fLqHuRWB/1nZE31KZgBCg+pJGtb3P
peZ/XYp/ngAU5kfVjRkacdlyQCLaLXMEjD7rp3oU+S+fx6shX/aJdhIFjj87UlXWrqx5FWvyAx7h
OBeJCNfxAcBJmF8gViGpf6M4AmoNhA7rSibsSlvnhiqnY+EPirxm3mUW5t5H/c8HVRIzB2tOLdKL
6dXT/K86ktNVspmBztfwfDRk6it8VjRiQ+H6ndlcdjcqVWRURorerEFEUdCuxNO0Jwbe8MGCdiYu
U/EPerqihuxrjCp4Ir+x3tN6O/gXiHkymos+L5uc/ABM4o6wztrytS0UufxThEujt1l+nu9j308E
/UxQtuki+6EsqCNbjMRJclWf7028XuXTp3RuYCUhNUD0depSrnIdme4fCqQfv3TNh6Fu5G3sMW2n
Sq1TJ3pevncK077PbZKMrOO9zhK6W3UY4ul/rEwYvZyu6ZFNGwP0OVooz4DTDiIxQbHha3K1O12M
yBszoBrPldq3a4iaQrLQ2mmTMGUwv5NtWMJZG0LbEjEUtggOOBa24cgpxM/LPmF7PIqywCWoZHeD
rLfhEqfTiEqqKnd0RJHwjNxne1yTKmosSWmEzrkUMYNHoIlVlCgmFWkbw20hLs7PuO/kons3PVR0
ZYNtKNHHi++GKztV3EvHqsTlKFgzgrG10pb1U794ZePLFLEMKKBn1yONJgHhnX2u2bA1euivKSQL
Ph9MxgCvBrnqAnMRvbcDVzJd+MYyc7LTCM12rKhVarhV8+zkQL/l3e0cqFQGSymbUubq2kBDwgR3
ywsuKh/WPmHHYThitvglYskYgjP1iGScwepRVHmNgSt7oSGDsYBT6nh+GnQ9eqoaivIOEET2UioH
PJOHz5BQFL+4sESt0HQ2wt4/seerEfZezYQD2Is44zu6OxcDwoWcaw3dg7bQgNWpJ3PScNy5y4f1
4N9ANMisNh5dtJ8BiDHCXTFFCaaIy0t5XABPFM2+65yhbFl5ROyflAEjOH4+7rgHaWBr4J7DxbuP
ggpzLe8LUYTTGb3O/Zrcptn4CeazpFq/y3OvRY7SiMGRewgFVitym9XFB+EeTZtIwB8p++NdQG10
MXf+OSze9aUleoqHmRuJthBeoLJxBWKpFYVRy7qLPLcdWS53Ro+oUrf1H5BEPYCBEhhoGJioILes
lMQXaMnSf5aQctjKV6biT2VR+vrSEFXVWi0PxtuEeNgtc+BZTLp+w5g3uVZ0xFZnbwFlvfj1W8CY
uCebkPwvpxvaXwQKnT1v4WI3yCffVYVHX7Vt2nLcG0uSy0fkxMz54M4E/lFP0zma3DNmwuQo5BkI
uP9LgEa+cPIqNpFVJpUFwAAOEJXSC0xa8yRLdKLRukGjEiy/YDYmROtetJZduubICH1anEZfF5pc
/Wa4a7RBF+udEa4degdBTCQdfsu6WfsBhkC894l4cPOBcXkEei6HMdPVCjaw7ClQoq2JOeYDb87m
ClOv770O99jvY5GOO6+kyfJJCtlMSmVp8c5FwFIbQoJHueDkj15tmHGgASxt4iGNQ6Fq8HyzBw73
otq/GWaZYGYnkSKVCFDwIhGcKKTyOZhlXfGSDo6+MQPiHbzKn1b8yWeaNk3/pib5qde2QLk31oat
BSZ3uOIsc4GwapKudw9DYpeuWWJWt9rVR2RavYZtQZExu47wO9d5SDu9QNSUBnvTYqVHtmdoPPn+
766Nyy7wUMJZzv9zAjm5wgR4XWxnZ+YPUFJAiaB1D4xIUFERYHCaXz0mmHcKUEInfG0io+gAaD9A
7XetCOH9l1c1jWKyygZMNQ8YToCdeWE5U2AD/srWsCmQByaKhKifvMNX+Bc7kP1FCIxpN0z4Am+R
Lue2cu6/ppxJLJ7Oeo68+vZmKjZXl3PNkE2xcxnPZyix1TjwZZOZn9u5TEl7VK3QGo4jvVgLp8QX
wF1G33wQuAHdTaP4ZqkweKUb6nS+s/NhjWnpQHrSdGAMpymTn1YzJXxyazqX4jKRiVX4hjCP9iT7
12Rp8Xr0QJs12c1JpMlof4fbE6zLhGwraSvTRazcv/xhB/lEUJfJt1j58d8GYiw0P3TGrzuaxRXe
aG2iekBVPULvcga3WfxBJYG96Kc9h0NHJ4zxh+OZhE2frmKqBAT/x3JDuHdwMT/MkrUtLMR6HJGo
quj2a3Cw3XlaSjNomZenYUFJUOxdMw0SA9WbAfm4dqS4Dp5zK2eX2uxRFZFy8wScT9qbAoqNupcm
uCYki8uXzixk3J/LHLrOol9qmxjj2ApTUPqKU1KY9E1EsSi41ZNcAzsb+j3dWdU+ZTRvn1ekijFu
dHxU2kK9v5EIhehyM36abbegg6+Giw9oXbZ/8RedIh8NwfD7/+4tuCyvKBc0q57tj8aS3VomCwKP
3qZsfhsEiF6lFyq5oU7lLEodHuE7bUF/iw5jDfwIYMyFTh3HDyl7dEGx8hVh+YEEaLH/ZoTOwtoC
P8ammVwTgKQ0HYUNzrooWDVm4Rnh0ankwijurAla7VsaM3SShkY9Bq57mcBgiC60rGVFBmXeGODH
1ZYDDSR6ysqqNBnFhqD/gmUFnjY+SO6rQdGaPgmoDbdBCB8zWyqKtZoVLpFlkLd6gR/vBjEIhyim
5NO7tst+XjpWt9wWS7erQwnU3UbeMMudbmBf5Oe4OzZaE8Q/c2phA/cPwo42gElFlezcPB5O7+g3
CqN1fiUxRuWrHEHtD/18KpftMoGMJitEX3YqPZbIUCSJSBLrny77YkbSJJ20QnF6JNqvQqpsp0wu
VzJqBKZbYZjaXvrA4/ya2XivS9eQS3rq2hKY6ueRJJZIZ9fati6AbrDNrcKSKth3tP8yBbkxPKNT
V1dS+amJm/g0TbRRGhjSbnI4bIHeQZ1pDthlDu5MwvsI4fZAoQvy8zNl6RSXZ+Dg7hqENEekWN19
LdFSqo7Lr0nCr5qmvBseaNu90DwTObpuk7qHp5P4G3Lh/kG1TAkrYIuLwjthuvV2weitDW/wNWQL
gnuidkpMMs5rK1J8WX0tIPP+R+LdDk0HR5A/3qtL8HnANgBUKYHflyCHoiIYQYZ7UmHqQaClvnkX
T7rprUO+GpKL3UBxkczIyGVsy49ilmVNhNEKSZI3S+rdwXGbbz9qM49rOvS06el+ClQGV8gJHDEp
9vcPhkFhdDHFJyj+Wv/k79Tt6W3YFKwaSWHmJXNZaaA8yfJm05hf2vuzXvjr7VSXYwc78AgQNyb5
KP3tdg9R36ya8HavXzKakFnWxWIVbyTO3hxdbsXHP9qYd7TpkAVBLFUXTSvzLyE2CCOa1fNUHoZY
nqVW7Uz0ZP4SQkUuEyeDKh1MpRFq6l9oz08kk0+JxiFNuOiBbsqJ56vTSxsJPpkP3JJqHqtPC7SY
gXMKHD8Ad3ljue4Ce14OIOnLDflBL7L9/0JkIeZWv+0AJ89aiGUHgMpoCwvRgwUzl54vl+pt+WzI
wmkSpj0nlDNYye9tYECpaXUHAkkZhKPVh2oC2o6O0DOWp7p/w2gwylwEU/wjgOE84hjakWSJpKui
fKhVzN5USfo3tNeEiJVM7UO2OEkrYCHTAzwlGrax6x9MD9Mnrd67lo2563hms71wo4uA22Rig4nG
XyVAxWszookr85FJJ78y1Z3GMM3KOsSGm/N0wRgctPRVHKZ6kEx2JlInp2gfHANwlwdoMvrtNcD0
1xpd8Wm4aASFOQesgBEgU/t1u1y6qIXJS0IqTKrYVs3J4Ld40L5C/TnZdfkYTAHDZnx0X2jPNPu7
iMWWuzvt+zpR5jPGINA6aGZ/J75vqYaDsChnTOBI9yVKtqF47UqbKqPgE1YvfKxzg8OIxW2ZDVI/
dzUvL8K5wHKeUKR75MBjQqSeG5mS5Q1wWgSRbMXQkYvqVDV6x0+O+Sh8KXQ+QCYnL36x/Sa//OFR
pYHTZhFgdAJq7Xd878al3XfMYTwB4LuRlO2gFy5cywa7CNb1cjyo8On0UQ5LAMQQRBnE2R/ANfHz
zI4cjJn7hzW6CA5GZXjbtdIPlDA3mXPu+TL2Xu/y9xCWXt3VfcsKyn2kEf0t4BYpWOwkwCse7Zbi
U7S8rOt+Wtpt/1NIa8sz19/Hf+eX+6hSq0bByPM6B+BITaT34cB4BUH0uuX130yk0WQwrPbgLMYG
bGtIhGR9oYmgQfgkvtbAhg3PPCrVfaY3+FRoVbEwzfMDyFa8C+GzF502qlhmq+bnVLkhHdGnZuC6
Lsg3oO/H8zYBXUzWS8loZsIKsYujZIwMlzICSTkJQgKyWsvdyp5qjFJ/V5kQh6wIw7jhq4L3mQkc
586a1ysGM+y5GTppFaVvRe9t+rmG0tI0MRxG6+OIufARcPni3Ien/apC8bZKgI+NFIpq+SsV6/si
QXShyfAl2g46BuSed3YA+gmnL5HyA8Nkn0/mYPkorleM31VsYAAVfDd5hAlis4yQRmO2kfMIejsn
03RS4RjxsR6kGctV7S9mqgzs9ZzZPNfEzguiFHiG7/RmTt8ovsfquXfoORP+ek/xgp+OhU7Ks85N
351GMTnKfjypQE4gODurDJJ/P9icexWuvfkuFGyVlhwTVZPh60fYXl/+drqbmSogg+9KBE3A73IE
jkCKIUOka+A2CkcSIrhm+pcAThbqnKodwAhvt2bGyYQqIKvBhZ5V2F2MjQ9UyvKxZaE4l43M7fAF
xO/EiYwi6Mcmx/WWsWDzYWJdYsuMl01hUzz31u++DlEV9phlz7+DRbSw20/0QjUSrJYe0zmd4zsJ
kA6uHpEir5svQuCEIvx01Wkdwy0YIbqIT9lyjc/oyR2seZLWB6vAOX9qaYw7x1XipRIf/vlKj6zb
oaRSiv/s1CMepqkrGRRnwWeW+9fju+7ahp7fXk93Hag1632SovOcdupDu1MW97iA7PS3MPJ0wp76
viZMjO6gZ8DArJziKkcrT3nyrq/jEFs/vuygYjLn4iR+M2OIbh1UVtPYETlFOEwgfpD9ummxEy+s
udTezU50XNk1l5slFG4r1Ix1CWfm55klmMSW2SEnP4oZh7RO23rNEyFJpu9pYfivRxuFm1VVyD6S
cLvefC/zO4xDtMozTiiPLVWeUdfY7ocFrxNXbATAxLyqjaRRERZrIn2WOAdDxUWUYWkbW022IGmY
qV7Cnp/Mcoz7dRC47Hk1cgJeZ3//Iv9gsgi0h0Bk+fh+qtxY0dGcsiZiNet0irOTdfKOh3AMvSdO
rvcy88b/v8bqSp22XzdphVg3uS8WIdK+snElJoFpiP30L5Nnia1Zoj+zKsRMh8tt77q4+AGBb8UT
QpUoxqyAV7ngsu8V5wlxQx4TKLd/Skvh62UnYefNpPJQ9Wx8gyFMApNWxNPf3knW0UvYa0zdLCry
DEn2W5+sgUt2KUWn8sOteiohoIGgsKGe6tGKqVdc8SfKex+7H6yo4H5/oId4DwzJk7Gw3JZn3110
xXwL1rgVNs7FCU557U0ScqHLj+y3ukH7MTGo1ZY/4TymGViJebGPZl7rTJtF0HLAvQPoq0bPx+L1
fhqkj6N9eTPrnfOs9aD+0UGWagN5WTkkFF8EdIURKrvtD2k84jl6E+dlreOnlSuoPKyHGndQCT33
OCRRO70dH37gqK3G47h68oKsRgjHUIS4pHkKmJ4cChjV18wpoFayk4d7HN/4GMesK209Zg+v+Nit
KS9T9muPKWra0iJAgzcUuwVFyYHhC7xq6a601UHqZJNHOwOC64SrAWmUHAC9PyexxsrUMBkpB3eU
4S/536koxcMmCwutoM0ipL/n1+fdHORJ0FUIl84Vd5oq4C+WzPhZveF/8w3Er0DIDYXGN0t8Fnhf
puKplRgXfpzyVne+Hv2Gypb+bQNDchbIYQ6apHpVOXBgSxeAie3D2PQcNImLlAyP7GPsKq0ebN8X
W7HZaVX2xGR8LneWlMfAvTKBOf3wGk6Ayt4pXoKVnyKZX2KamGKQ20GAY+5d0Dq1h3chy2wDfjuw
sh71pthjonA+yc8y1EOoWUCGJ+2JuTwyyNXPTBr3lgxuV86KoHtJA43ITFXyfxvW9+vqctJ8mXuh
sLHLen4US+DmApPAqDj6O3PJfK55PI6dFTrzHAqnr7/FnYxOGgNPBeq7GMVy5Qol4NB1nxaHlejj
E1YHLLPglhgmN9PPqkep+x2cER6qYk6NEaiNhqZmzzBOiasFKTU0I33cDYdzNFoebHcrQ3CGkHFa
ECoIkaWiAcZDvKXiBVl02tWOj/wJwNCL4nYfY8p7vXIq0OS9ga1MIrGv/81/ovmduFCIjZQuXNM8
ZVp69P0jUlyx+1mAuan3AxwS+sZ1PpxV1pDLP5Nv80FCgihbDLoaNeNx0uNpjNKCPJJNEGCWZ9kG
K7QIVdxHGfieSOcNwjDM3L+GqQrgXRYdURcHzW5Y1Go7xEG+h/4bWiODrHB8uvtovx/zFk8au4BR
xXEHqdUEFRBJmy7fCgkYUhu3n+rDHpdl+QproPHrPqHHckKjj0mPsDmRJDfYHJXihPuKviskUCnp
37DC0j5GoYkB6BaL9d/KMzepQR+Uo42mEE0b1S+VtOV19ncFolCUzX8HZ7w/dNNG36EH6LW0LYhc
4nAK4UybYhXkNUydbUkKAP6aXPFHwC+8BJWJRPwS311anIq4GHjVGMf+BfRsWB+oyxZnwsvI6AnZ
kTRVIrTpOMAq20Dqy8iv3/4RFuFSs9JzZbHpokq9DUTlsOqQTYo7u/hF18F0dtY55rluyWXDPE4Z
gLEaIwmBUvIh/SX/OFOBoujwdNma+DfSEDTEgC60I2FN3ooYUnqTtvnlowhBxUmblhuV7ufKuY22
gLQwpLjpggXiyVBHs6grMlhxepO+VZOrMUkxg9ADvnbzZi+BbauZzJoggeshABEPQ7mpeX8c/Uoa
xNVa9P3VmFKgGkhWRrgyY/RJD0ym3HCnS2j7QlUm+aQl0usFQXGQny6ZiIZKcAndRgCl/Kc5RXAz
2SnRvogpyj1Ze6tMfEa9QYpBec1+KJ3gOiLwCxUDQf5r1JWcBgpd80Y2ndtUvYuhTWP+9H89r/fq
avpDAfm9IfbjjQD5FsirniV3baWqiqqiuigsonbvfPuoWVntIHGXI2uj8lcBn9mGs6wYT8HectVg
Ydc+H2nqwiCYeF8UOWtvUuamR1GGzYitCwp4LtT0lCUKi8tMI+qJFJ8BVR6fEDABJJV8vZSTKzBN
rtUOAyiPnM2HQX1EvbEIU5DfNSgsAiIF6A4HC95+0L96lSCbxwsw4IB+PXOycEEezjY7b8Mr0C33
aGTBdarJPR3Fj9Au5PVlwhlw6jnZiRqZaxY66Nqf9NPovcQNvF+8ORRCC3ZsXdCSDPwCaIqysXbQ
XoklhxPHvWYX065wdXb2exqMi3Hxi6oJJpA7qhqruxtwaWuabsj9JDWl2JK49chWsy8ieZiV+nxh
7RTT0vA1KVGAqZELWzC6lrpTvrgLhwWt+WeLr6MKbjSjvv4KRceXewHqND74wKrsCkLb11S6HxyJ
fuc2NyPFnTl+f7FMAhvGzjldveXE6VtazKOskl27YZbQw+lOoJ+Xvkh3XPzm2iqOAB6RbslKhwuK
TQx2HZRs6hqKnNg3NrD2vE4CH+srkZBRzQOIbTHz0O2YnPY5B5LEVPuD198b6KexQo4iSJwhswbW
tSeTMxRU1KaMEEfBo21c0XH41MjVo+v5UPwe3LCDe69SWrwtAoWjxxwAxjS9bhd6DDkBkkk2Qj2x
/WDlk2uUcaRcskq4Ynh53RnFwkdxaNLdkvOTZ3ciJSISrRbLE9qdMqdW/7EvKBhggJF4hGCAV6Ik
abyt2hYCucl5MC/mi+eoTakQ2yYUVjMfXm6ZEpwQ3j+kCJ56ogeszXVkOwNGvxKO1i+fNc5uKmwy
cotJ9j5dHeRRk4COoB/lcd0ZnrTQyvdjmjfJQr2ot7V1jIyrpfEzGKwA5N0KcU6N+ScyLWhEw5Go
e+p6+xEVfx0b1J0EkZpn26HtjdMg6VaAk6+PHjXKr4eC0awu/nQbPChkKllJ2tguPI4z78Ex2sPT
u/BvMBQmDfGYuy4xWGb8pp7kXYgzDr88dRHV0Fs+IKdZPII2YR0ET/kB0CW/WRIL+yaZ6Lecdvk4
LpD9KUW+Kg1BGyJJzMoQ1c9hzEGZg/qrcE9XILxvGuZS/Z5aiT9on9RzMUc3moHowGBHkkyAmo81
snWoMfqVvcEo/wbzF0ayudIhQQNN2Wri6PtWDHoJFd1am4fScjgjukWFkZbb3AnBgtkgvGfppVZY
Z4v8xnkJC/nGrItuHoSxDZX/muF6huKYaxjXvzkJ4sAKpG3AgdxudOcioW04ba8kK2km16OQblnP
mhxFl01u3mJGVfwvMDFkrLgs7QZftkvjFLxQF7w+XRcaxRL+RUByYsSYBLBht+2JZ0TCpvu0PBuM
Fc3ggs4M2DPSjwpV4x9/Hd3zEdw8tw/RUcQCclwtFpvf8N7Sayi8V3+pRN6m8sh5okkwwgkBtlec
AjwHlaeaZZtjicJYGNA51rNNR+DDysWWgytlkYTRS3H6zR/5Djwuf9LJfSc9y94VmoExS9KJVLd2
EIi/S3Oxz3PqlevS6bs+BkvtEv3JdBvN+relHMoHYSkYEwHw+vaZhUPgyMhA/HXFWhjsf11TU/Mk
encDU2bNSxCWHkQ3YfCI4FfBFV9wZOZldc0/fijaVG0QaSNtHyMIoFtt1A++KIKm1Oe5JoP5z0BO
idtKuxFYMo1C1/8atFLupMq7trczIQNN7LcsILCKNHYzwO2YNMD9wTOAqqiAVuNtVn2VGH5k+8Qq
RzObRD5wBrmHNGU3MoJzEA1DofCkwPbfZUJWCVdbh+pp2n5crA0Y+1aFubx2M7rN1PfXvYMLRtxO
ChwE3eZYSsSoieBoccRPwYRfvdulS20tHHXimhMC+ySZeraX+lHvKccfOR0HiSa19woBr20e7nZ3
VLv7Dlunm32nect1y0TrH0iF2+CP527nTfmacaOpjosjLJz/OLjwo7nYgWf/1rZpGFA+IfQI5gIa
JAaSdlk5s358YxWo16vXa45M4zjmTIhsEbNXK40HnspUf33ZJJX7hgpiZCQROAxeB3v1BbDSduBN
Nv4DFIxiMw6ak0w7N3OQ178STamI6gVgUJGL6rOAFQwyY7GDCtxUhFbow/ABoqikVctWT0LeBQYN
sysGXOv4fW5T4nj7FdVSLz78D0xR0uNrxPcSkgtL/R7QCHRLta0KAMhCbnNUIFWWEuLy711h6nuU
s4xq+zEeZ8F0bvhVmhrc9rhXMVvH7/IQTnJLrafclXhwQ855ua6RSjmFfHZ0nbjFWTFlaQ8GV8kn
5u6C1pP1BPwdfzl15c/68pynJED++BNQ6TyVS4ruVS68EJy8rKabcIVhNFGgw7tMgmTIAhmlScw9
D8CA7FQKjj0GP/pSKt20FXJIKRfVNGQDtVv1geAKcaavTVTczTM0QZ31X45D1uM5uL5Tf103OXfu
NE+KFrhUfw7AVuQZoisAwlOnMPSic8v9sNyxnakdoxwdttmrGaQqe23JRNjStE0oD5DzKPmdf8qh
AsRWSSRF744TspqlDmDaaT6uj1LU3E8/H08+gYjGueFO3ibcmv2C+IvmIVhONQrj0jlB8aB+5bT1
n+Z7Jzc5qLIQFfdEU5VyHTcRRuGGA+5JSkGpFW+VFOs/l36nj8HcXkEMq3GoWjDLe1GOUVhhcuUD
ctbvPH8IQVeagqB0kdjlyLRg4UlKJzkb5aGuNQnliDOtFgyctn0UuEfJxeq8T8nkOBpiFJTXZ1bv
sKyEp+Nn+UuTbvz7l+B9AHffhsACD8FPTIHXUB2yKZKnpuhlrOZoEIMF3PxtLSZpQm/b1NP3LR2l
yySuvjdzYplkpL5TPfSjzqyRbHrVkebpJJ6hFirDl02eUdecEIM7hO0hsCoonj5QP+Sxwn1uI5KY
ewIjDH7hKJx9z9pV4dm7HDBIhr+rQ3/nzWGHuhLhnj3xVaNgy4E3L1h38Bam2lYbvC5jYJnQAs3O
3LbU1VKzc/r5FKqayiyM3cRP8FI9XNv5C4vpycwbiINxBotzifQDbt290uaaNOSkItw5fqDLN/nd
mKyI3JSi7nAxZuJBuBNGkmhPYFj2uZ1E5BYHJHn4NjAVwGaiPoHcf19ZjiIwMqnE8+UR2sL/mYKQ
gw7zRjhMDz4nYEujcI1jPnMqsUAGxwOpYdOSn+Qj0FitLn/FjrqhPP6nE7Shkedsnz/wPV6WUvuX
qWOarR+8KDh5Q/BWwZn5Qb3Yfdz/nsbp+n1eczecKDQVviKXIlN27WqyKg1/C39T6zxyh73Odl+o
ocLE7rWM7+wkqxRgDAdsEwdKfDDylLV0Ai4n6zNHo5XAS1ja2RXuEid55Ds7ZV/0zOa9n3kHxGzd
D0bK37Rt5An0rmw9pffe43vvt/hDvkrpTAG7tAsrpCNW4SZgr1ZAwaueJ+t+EwNWMCZoQit7kSUQ
B3l62zrvT4B+tCK4hN4rgYVXWoi3cdk+UZLLLSwsBaWAtVhrrMVjF3CJ5gzbbYihMibzwog4blHD
Xj4Ei/CNlKk4TzLcIiHcLtz3sZYWpzofYbWBTt0N+uUyIRXOQJFhZBzXRXqx1rzv48PCJuz845Ic
NtVtt28Ot/iWpEmaElpWA4HOr8tpTSrkshdFhLoLMKMTKaHuh9CLmO15Xso0XxFlHqHelpr9+4eH
n32sEw7H4axEoiRNY7jkTtbXkriHZQpx9DOuRrG449XAtxAh+offNgKoZSGrxaLbyVHt+iLEDe/0
4bYG0WwjHIUoFyyKJDQwuUnw+UBOSej2QBf9yXDxJijaeVAt5VruiKgyqoXnGauYhsgjV66/csoB
yXN6Shvi8Eg9szsnDlkOled9yfD8+u/74Onk1aVA09q8ABEp6zwzVsehEwSGRPy+pMcB0b+th6VK
3AHvsxFZthHDQ9lg/J+73u+039h7XU9y0XO4zs5q/8JPVPEfiH77eOV2J50gY4MzaVf3uu3ZZNGZ
q0L2CFDH5Yax77jeClTBWS2pn83G4cYiJr/bK2fJmSiI42phTJqWOjnt6Tt2rE4gcQVtlLYjWz6a
glIpLX69pPEBbUNJo7p23xTSN91W0EMlSyfocE7O1iHUgXCoR1vRrQNILL1zH4YgngZe7P0x+/1C
7MQY1XlrAwBwfHZV8wxElmXJzV1RtIQXc+LiMQGlzwaCc6WsYnikj9PkcKBRFQZ+ZtdfrZHmpip7
AfC2rvzcscLI15qInavjH7fOq3038JtIvcN7JOpEK6RMtxd7+VQb1KtJk009VKuJoecKl+tkdAFx
KWluLUhAXP1Ii0YaQGQ/5yAX3fOSEljSxrVDAFWGbFYljnZcv3wBjrdMIUmu2In888PntSbQsB+4
g4SWjplNHlkLeS4vouv9smE627f3RC8+wClG3d4e1Ib0U4jEHE/+mauJL5wwfpbl7yusM2R1AleH
GxT7W2H4Jr9cg7gcqTyA6MfLOEyTfmMCUGr3b5BYC5sA4dfMWSytoF8uJNPLrEvsXB9i70lDvbcJ
rVbtQ2Eh7V1r9TnvARw8Qo/lCgS5JV5Sj2uV3PhYfwTD6tkLBxyY5ecuwND1lylkDZ3XUWJXqPhf
i0e86gY3CtsLxyCTmF6gCTo3LfY1WDj2gny8y3pXgleqPvWumunFF0rGxf2maTDbQgVlTnKZIdje
3kXZoazgYP4CJ3Ecqqc9fkla9kvZLhyvqkou6FUORBIoEXui4VohwkePJeO+QYdHcnzMW5rpl2Jh
uOVBapKzwMoAUmUFHM9YFEaRafUU5TS9u7/hfG6ptGEJ2CF6JQiGYkN+VnijZkdIjOuR31v23g2J
Dlc5IhBZiWNvnuEdxU8OVH6xM6o7hv54XSKhMVikfc5bmD7vzzG+njrqxhVI2amnPOgv8tpzE1mv
DY/1NGJtmSnMZ1rgqP41Eyt2J9gkzlUwekC9fYSzqfrCbqAieb+b2pX7FFAYS1EWUwrMv0cu2Bbm
BzAY55Ib2aTcS4y3BLakeQRInQ6ZYa08Pfv83bWmkOjaWrd0aJlignjEy2qDZLBSkG0S8Kr6eYTV
gwpbLOIfSTL/Ku+QPwHso72wTKJbwfFi1JqY3s1mez9MQ+j+1RA65be5Uy88T3rFYTvdbD2fpVNx
ZYrQhJsAxBXTvD3f3HVgv9Go4yaV+ejUzI+f7q4naEfcfg3QaGrMQAREPxbfPjkvOjeuVax2JXv6
qBdnTzN2cWQAZpYzk97g1OM0WZGFbRpi3eNRTDWmtZ8IVKPj1NZwOvAezJQRtds7SYF39snlapmZ
jobsIAclTg8hk3yHuQGyXZV+FUa2lgYAO0lU20730deHIEVaztY1J5HHKjHbggStVj8sKWGxJJiU
w+5C8XEeI+iJRqjyGzZiy0DAcic0RouhDHlVjp7uNvMhX+g7jzNuxluvPqk5VNOwXMsbvnjXq8ct
bO8jwkpdAm6roD+dnyPFVBel49xHgIa/6PXveqMkkW8Nd3WYRIzH0/gX+63KYY48FELAHH148sKE
rkZwbLmJwoam1vCtj76EfP58yhETVQ571gVb+PEd8qIkVtxaW9LkZHeTDgcyAtOFehVTYOodavR3
Tlyvjc+HyhiDF6BtnR0h/Hn8Q5AHDwwcrAA5dGE7TSS2/2wYaqibIrHBjjj8dtdtpioZC6j+G4kH
W3hTSzpjn3ZZ3X49F+4lGfqQwz7kMjAq/Zsx/JBWF5+lywKHi9aSDkNEdndNbI1mQxwnCeWijalT
aTWMMr3JYXeUNJl4fDVAWlx1i03VTwLd5ILlse6ewwkOghEaTYRwvIp3m8GWtggIQNhdZSTnCiyR
wEBoZhC3N5gKEuOiFZSM+vD/hwDGqgfd3XSQsM1ikz42OT7yu6cr5E1zuNLWAyF4h4o4/Omjrzo5
qkch7ulUIjocJXqbaTwHnuKsOKCEUe5oHtCJLYrDRFSx2oSsVdVULQ/5yBDFtbMLhaXb9vx+vb5M
ho+eIWx66yD3VYyiIYjVpNtjBiUqlFqpcVH3jGVWQVNOkvhcK7MOcM+ZcE/kO2bgHKn0+CzODCHs
SnDIwhYB+8lXr3lLTQjM0m0r/U3CWVQm6rAl0MerewuxlWX4dRDXCpQjWdCL3seMEU9wGJJc3ywr
EUTDYi1o9KwGKCzEWEKNQZUuUubX0ZfcCLJgfUCywNWMe7QOHvSNBaTntU1yQqqctCP0+Ya176sk
PX4F/M3oiP/BA9mOcDvr5nIvLeUi580gjUzzpWfcP8uX33fpBS2MhcHFwvosRDL6xTXGof5pexd1
EhwWzomXPNKP3hiVn0Y/WwaOl5YlmEyDmtkzGXl1ddWJnx1JOd/xVFsVWKsfF4IWenD5y5+v9hbx
kl29e1M4aXEEKIeOwv6k7c51gggFzK/itZq/Blw1HdYDJiiJWpdtZPCuZ/GAiGCeYs6FYA2CuGjg
36HGNWVRcwBQ6o/GdIX6HBnzyEmMNfXoXKd6NaG2/DDLvW82c8tdi6VAmft9Fo/66W0PSNKiyL/V
OErgQHhDspvhl6I8xALxHnZ/7i6SALRAyhe2Jis62BScgUJoUuHLVxjdb7qzF6Qt1dLzVMiDRIQ/
NPT1afBeTpNagonShlnAuFcAsQpJO2/Ig61zAyD2GX81uaaislUHzDZKi8Zy+n2aH13wBjK8BQaB
yFKBTtzf0rL+2m3HEovFvOWgP9AtY8z0kMdtFuXRuDOLCAWqY1nnkzE8XW0j1nlafLfimO0DQ2SF
DKYdjiq+ANxSDqoMq7z4bNxn/Lu3OlhPWSvllLYk/MH0KXiMsE8iXMtKRAdcAtBoOGbVt8BtiNKH
ts59R9pzMFpZuocmL/zfCD5B3KdiUTDb3AjjjKfuiqZzN/+Sa2wC64Do/YEeNv3ByH4/a8cCpkhl
3ruu+HLlgFTG9VaBRdAt19sTur3uJ+zjj4u0raUtCewPk0z4yMrEoAepEknurWDWM0vKbNlHD1gp
jg8b7/+Kp4n1VG5biLNMwPAPqm6cJa/6WocsfXj5Yj7Yw39RCldEWfkOtQgIcm9Rjvq02gWnxd2Z
bhgYqMRP358l2pjZ8fG3mutuGNJX7t1fAI8iJVrFHSRmuhtFaRS9gxBJK6hLFkav3kxCa29K87Rz
jb815nwfCpcSHt9huiUFn4BbEo2UC6GPb01X2UnWTTMV1Gjya8DvoCr2A8QDvU0yCuLxr8EuCXTF
Y4EIZJ87L4NtWpHDXaGRPxqq/8I/ldl0F96ZfaEtP/MQkHHSPtzG+o8cIp556ZR/vN92l9sIoA1e
gWcS4xSl01WYRKYhfVAHPEvotLFi9CSVKth1f9BCjwqHmqM+LO8NLYBskzfFqUNXEbXPgq37n32Y
SKdYTv/T3fqv8NWM1LxmvSi9+uebrVJ8cgPrruNMQk0JjPUWEc30qerKpyhkaiS94Qu9em4c9qs8
nx1WYs6+l1JBeo7KpAZlGaR9AXiM5J+gBMFQLkbvk8HU6HbrbySyHsGJug0IrH4HD8oSCyTE/qnc
PJJazQOjQu4YzajdV9a3wuGFR9I7dkvr4BWZOyEISvnKh0sTjRTb+amQEEmvRibHDPkUJHxXaLkQ
fnG9Z5hPqPUPo27Zw+XyNrA9lKHG9LdFeAcL/MEjk0MXBz1Lw9JUAXzK6s1MEE3SgHjonDjAAS0A
PdZUKyndiXs5CdPgwvU0SV5FQeaBLZloe66B7d0b/CEF7l8aWrUTpYFgYfoe3WDtsjH9wTzZ7fZs
R0G76qobtfSGQsBqsaF/2Ga5T1isSKcXOaOER8CL/qrA2Y2tB1SA9KB/wjOQu6Bw9JU5FsWMx/UE
Tv+rT9GksE4ApuyKej0NIobOoadf/v3efw2GvmY9VHAwF6yR8u/W1nvOwhOI3AU4A5kV1dNkidA5
Z1PkEQcM7cIhieK0q5/YgcHHKs6+zjVtZG7udsPmBmI0YSgkrxCTFtnqIvGzhrTIQzxntyZohnYg
2sKHdsCEo6IEdzkpemvqsr7mAeOXCiDQ3wtxIAaf4cSXVou+Zd52HTd3IUI9JykR+VJEmQtdQL2G
IfzJk/tm/AyWRzaKrw7v/4pN8KSZCU+1ydRvO094eKCatmVS3KFzx9Fxg7Fiul7534kseOj08Z+L
sOU2M1kcylZsh9dCiu4iV9sHxFJy9Xtz10+yEWzJq4NwWbnxpidhzozZixmvz77u87Kn2YPaY3no
iuMPzbOaUmDJVSrezY/viMwZh6+sONyl181J2TWAypcdFnMiLaRGZoGfDq5r1OfJCjR23c3naJ2W
Uq+vWAGGobbcfP8cWbUf9pkx6DpbYWpVcw7w/IspVe+gVbF7kDn1Ltr3oD8qZC7+u3Ab7hzsv8LX
+h848gG7dVI7X1QWOmwUeY98Ado78zHYbiCGkpCwqUrgIvggggcmnBP7K/EvDj5avkcReWzyDMiA
oNS9ofGhMRq72L2wMK6cCgPZgx3fQlR67ADZHYb9p777u7cJLVA1q5CZWq2We+bemdq8dzyi/trX
RDo7R72JFKWGGy7JhIZWNtR16JKok3LZUi1VroEqiWBCpda1dTzvE6X23s1+uIBTDHCYY1Y+npxE
IHkIuYc+fz6x7Xrw/bu7gID/7vfM5qP6Hn0shGNWts67eBf+bIs4xFzpJBydl+5oKiIkN7T7Y5uv
UoSpFkXHzphwcwwrF0yMsRDgRXAm8afkKXlEZkhS+Zz8M72E6pVlWJ57TtQzdUGHXpkzqUbQUCsX
ADunYtfdlSyuJCq4s87cummpmmUarUwhTlgwChx5jnLOAWO7QUN7RkJlSH2//PS5kRt6JazI4DLM
nIjI/IgjiAOz3GQlbPQwIWZPMzGvPK/sIfRd7c1uwmOZg5Iur0eBMzQzus+RYKucNitXoGd8mqT8
Qy5e5aGfcdQAuiFd+ah6QKqf4mNVCamWrDWiEaP4Y/ks65CBDkLEbGL+8462/jMi4tcypdWki3I8
uag2sT9fIQMOG/ZdapBRKxQkMWqTDmX/DIyxfC8R+tki/cCKPN9H4hTGBWdPeU4fTUT6o6zkCSkn
sliFDGT87DUxBjbZRXWj/f7jQRpjOV2Yixmm61Zy+DhAED3SxFZNzSvf9N/l0iZKW/dY1kWpwhLM
W9375X5VVdS4HFUCJXPtCGUbgoAU49VO9jgD5WjpSij20q3tXjLSLdMFSPLBSAOIvEUDtPI1oxSR
lpADwo8HfKt5h47wBoxKdw8Vch2gOGWK6UKX3K0dIJggdf73L6y9FRkHMEhohKQG4fxQEIE6Losj
23ndWPookKsKFpY70ocJiXIwRH6hxoIQtmR/u4GxauuZpJ1j+Q0dWl6zHuHkbEvJweIS7ARGw3+c
jEcUp3uVVwh7TtZNJo2rtZSdpcXxTp9mwUzF9cwf1XhUK4YwjTiAdnaOFlhEEuwg5l6mRVMI1ugj
Wt0ROvyeTyWVfu7nDN0aPU0/D5sALOeAwChs5p2PD1N1RXZ9fTKisfy9BVNlAzQ72knWXWmUs4BW
hZFrTIDgmUTPrV4iyvvjYnYIiCHh1RltIpiB6uP1K/M4B9fL6/kzTUjf3CV174P+357JQZhskexR
VBOpseRhiMj/vaMZj+5h5OiOZrGW/TlO5+be+zlKMr5IdLgZc771lhXA9c9m4+R1MBjzNBpxJ5Kh
K53nvC7H7l1VbwXnauZanB2QlNqM24UjhFYpH2L+OE27n4nsFFt8vaSGTwBdGdMLPZb9F+AMiUhI
jmhG5qIVYFCvGsgB/JG14VqhLAHdf/PtWaDlDXCXEk4DlA9FltbXVQk4CTMa5kHXkXpHIIQO8Ghl
OTMHQdkpWpTqweshIdyVgwSyPhtpGd24kxlAXcIKFzcGCaeNXwL/AO3a4W/6Xug8wc0GZr6lrmtR
Tahbj8P3na6IMJPtJtyjiXxlSgwiWwJ90a2FO48y+KbH6/ScTRU7hjb8seRR91EU/of52PGi5peF
YHL+0k6hk4hqP2wo1DKVgNy5kqUHWxCIWVvMTpB6F6tuzaqwgMQ4w/fIHsUOZJsh4lCJFaGv9esp
8m5lSkrkQ5hniK9F82neMm6IV+0gO8wHuh3kWjR/NGZXSLZCt3rCUjE62JYsXodxoE2UPMW/IXhO
AajCMYyrD5FRVD2AqEfwpd1F6ZKWJm/UMsAGZhG7SKc0dfVhM+4IYBtuxjrU+mfny0jpeY9Ul7ns
IQq9bMLHBxWMPtWS/hxUDyck/nFFCq6ixrWQtjtqViEKuNWJoMV8MN1f9r5gjRH2qFYn5mVePf4f
TsSs7MmOt0mtNbX1Rqxy167SFJXgtPNHH7Qx769Jx8mGMr8YqlRzqkElFklywoS8L3MPpCXNGsiH
wUMTu+hhEDkTkCI9Q4e7+vqXeFjtJCrHwKiz791MQ0WQOPp3fA3UMooBadZmm7fbTBD9+TY7A9+j
YELpdwbF5uF8s2SyVplMgsZuiOCKd34+dM8Tvjj1F+6+g7BXFR3M/WI3ac8ArMpJtJGeFELwv/Ym
jR9MF7sa7ecQp/+Sg5s5s4wPJ6Opr6HtldM7f1nva7V9Po6SuQmR46hNfW1cxVtIuqGWnEXAs/l/
kt4eP41wQpF5un61jIhGnplW8GmQXuukmFbXLUw906FaR0fPR6EoeO5hWecPZuwUwsVbuyQlV/Ko
ZFezmYRbD+usf/rn30dtf0+2pNwKR9CAgz1wXGMilkcvaKyP6hGF/wcvcAsbe3k4y7Emn4OsWony
aKNH0ev33eLx5DM7YkQhOLeFP5rlrn2qn8sRZp86qWKsr/zfsCCCvo9bPCrzFfGOHsrxJrMtN8bN
o28r7QITzwle7k/kiuh50wQd2t7ZtnUvqxYPzzgGKU7tTLyaADhOVcqZ1YNzPZ5FAs3QpXH3P0ai
Pj7AOX0FLXkn37NAr2XFr3rcbCtdaA/APPcYjwAgCUz0pD/lAHbwvh3cV1ZeknuAfEG62VU1ClXC
68tmAra6ky9bvn//lV22VhNm55lYkYW8vWLIrm5xvQsovGVfJgy094TGNzNjJXf9wsuZN03KR0jH
aVDWA05Rqn951zVUg9NULIEycjSuwGnd4aprU+tnrHw50NcuKFB77reo5U2ZXtB4e2DdsVQUEKXb
jhrqI00eRsKQjTfm1ptU5rJ6c7HfRhX5M7ynMkD1iA8iFeC9pcHyvRYLjHnL7RVz56aV1LzUG3kS
yjiXzsH6CdGlqojLcSTpZ/NSA17I4E31tdfXbBHPjXpyfeqaW2CJFNvm+Io/G/u+ZuP5H3DyR0Hk
w8oYOGsB5vjJfgqIvZDqVb2G6eTYUvZ/2tNIixetDm33xK1H2nbFFw6BKqgMDaOIsUrNNlvI0uQG
FDLFb6rAcF1E0Zy2BdDaMga7eC3GhTlulS3AjYjFl4wfNPdY1Cr/Buq3nqfZrJ4y6wB/4nqkDZBx
E32C+DTE8BCFwWXJeVKiTM+nyEmmlL3iW4JWANfd/3yBq10qEEZSF+zCd/dBm8cVa94Dcg4e8/dU
DMb/RtLGKZSjZbzY+GYAAn16VtXfGnIlW+gOZOArrMPo09D+zaM8mH9lWGqUMtOllGf3U8WzhxbY
duKf9t3MuFDNh4cADr8xAmzT3Yd187auxJ7B/rlRox584pq6UNY7VFBuEvBcYjB4dw+pdvFOjabC
6ySdF/eCR0aS0sr8rmC+lSHOHo7FwRw4NC8Z/HuDFNvuThU1ro4/OCAmnTKAf76QEoBTeORzL1Xw
g7cTJCTchjjVse7HPAGtAJeYt0jQwPTCz+KKZ078GEfPl7xsR9aGklR/tjpZWcolOqEyJue6Qbgf
Y4ciINMSBfugTsAMOn12wow5T8hrC2TSCHMpJ5SH7SSmIsOtT7uuQ3dgikKG8J2skE7XgN5kDJsf
2DjII1oiCo+iCaQ6bzbtzF2VF4jYR9B2qFIiv6JUtx5z/Om/xSN20DeuCpcjFJf3hfNQdyyqmuR+
BHmb8uKgxRzw32sUu/2BoHCwNZplY8Od7K83B2UY2TYJHKMM2ANIIWmutvaxe1694kzQi67AJmd2
VKElS0xYVKQ1lOKrJyp0+1aebbwz2n1pIRvAGlKNJ4P+IL/Pr2zciknuzsI8R5mTS6RR05WQAw6c
D8nhWLKJx61L0YUud5UEIIuxpM169BDUECZnChKnzgw3F/QnVZqYmo41QbJO7SlS3NLACz9AOV8N
xabFWdCDLQaDUiaudF2Op/QYCGjxnEXT8/mZeW+f/Bh+jv/yfDrs5Cdamguexada34IEAwsrjmIl
hLmtk9MRIGzySYhmKuz/PhSssqhNai29aIdOqCiiKE4TYUw/9LwFprc/9DEIdeTBhmSGCHbCH11J
6zn2E3rEsJT1ommV/cmSxq1VwC872EQa3FqrFvtayZ0laAusfusKSwtmpBY4Sg9GVtf3Ei1jI+hm
edGjhBwBO2G3MwNajOKHx6M7470I4pgkNfT1ineIAHBkRIZnGmsEfXqTEK2TWnKKOLdubjz0k42/
S6WH3HxEQyPYsKyWdplayrRJVpzaN1ZJUHXeGSAmyxJsRU7DEhPEL7J1h6DOG7Qm7jB8ltTtQZwX
lrJh8g9b/paJVBc1cj15YsRAJQkWIobxmJTyBb4wSmATnMVm0t6++MCNQ721z5qn7B8DmkYxlO8Q
Rrm00cVb9r2sstt62EOXOABKRPHG9PHlNr+JyIbygjgNf/xlQtMAZ27MFmTQM1xH4WtBCUpFsist
DZmsrrrLiV51Y2bYoX6p75KPLO8IHLMjcAZ/ESOewdwnwVIgnrw3HgjTgoBkqYX2nFXDWHpJRNsC
p+ksoO2d5sYeoKGZrMQTIJvOUOL8zN4Fnz15WgPi9b58FBl5+na/73rKQkgJIuGwwYVMhDZwLbOv
BOJM3zdaSxPgQIDkiDwViAKGrKbf6XhyAgoPXJNh+Dn7QfnbJ/yr1FpO+/UKaLJn9CyVlmL/KeF7
7HpYIea3rh9NC6tM+xR+B7L7pSkt+HfDmR5YHvUxkaT6Qt7FYHq6iPwE6nsv5fCyD6j4n1zRtvMJ
gbPDhXaDJAm1wq3Kegbdhn/eiULGt6wLs9KQwWfS2jbzETATbu4jL4HJmkyeyanRBWv6iWCyqqLk
jZZxUpQs1SqBQ3CL/GcZnLYrbtPzwwQ/UU4mZxUvlLcWxoFXJ69Rw/qXo/1ERNHXOmj2z2vSUb4M
J7XUKbXz4AcpH9O9XwQLvJ4KnTZf5SmnHMk3b/CO4ApfV8mho8Oqt6OJ/qNwp7lPQgogshhY+FWa
zl2JIQyCQrseyYRJzJy+XJAZ8SxH1O2epQAlBUenOtkvsUn8+MIzG2hpbUxnuPcMfr0ALXZthXvN
X0PzP/x1Df+1BipmRsI4OiV/Ls4xxjfNd8rOAxYq4rFmdwkVI1vUM9aAuu8Pauvpx5LMTkN2KNbM
fbLFxeqJpu36MhicMMDQwZc8ZMeRDm2JAHGfSFHPCmd3BmtbXr9sOpAr3qoz+oxmjqeHwkfUxSQ6
gTWn63YlqTlaw+4GLesF0gt6KfywD+4z/sK65b07AtMWekyCBXEBtj9u9vviBBFeERpmb6JZtAf3
ZRrGJCsP8kjMkafLcaWqe/LgffONOw3Z3oRiFYZIeb7BcWWR8sL3lo8NVR7esOqF6M1qmQF0JPW/
bsnGNmQBiB/ZOX19VR8bmTTvROudXjK+7e6hZ5CQHRQsJllu6YGAMTvXBb7MDKjEvnmYhq8CYoE6
djBqQxfutSIbaCIdq2oDbP5s2w2psSnGClqNPsqgD8rtSRk68ZvSwQIeaC9t6pjk6VSkp4eHJeWw
szH+1fc5JWt7dAnQVAwIteuDiC3RR06YcB6OOfwEeLnNXhiohK5WVRTjNKiBzEjI1KzZnFXKpE51
xup13zQ+7vwuz37UwKIoMGaRehfjZONZhWtBJpTkKSe3SxoAa2tNbfRs7T8Yc//DhEbDgamW29hx
QKwkVGl2duZbPDjJTPKXbqOVMMKm87IFo3cojq+VGNHR0fZnKroxMdXR3/k7Gm9xlRH+HOTfFojK
d92pZcInMN3xhLSVBumrbvwfBlxx+zciGEOsYl9F2i2P/YhdBlofdRD8gK/FIHLmHshCghdgmRs4
VTZiCnrKIvpcBNeTynVlu9pMtKclTpBX5RwRqHebieEhkVfDIU/saXMdQ90AHB/ofyuEyO12iloW
bJvR9ig30Z7eFQczgOWHo9BHLsM5mA7Zl4FfpA9V/aBsXdgVy1u43x/SqhEG7+hbqne3XkRddElB
HF5EQyYbrr/jv/n8w3yMEo9TKvs5x1cqrZSi7ecvUEB+R3LMoGZYK0/WgPqOIVjQVRJnghWOer9v
8j4n959utBejU712PqFTwAY7jqy2857cwUVtB3yc1YXYRcPPxDLAEbGRAbFoAGgO9KNP5u8lRqNi
9OkPCW54nCVx8Y43VA+OsSNS+zudK6N1s+aYRtT2T71Ha/4HfP0HA+Jcf9esZuTKL6RWaL4xLunk
LY791rITw+2pdQO8hndG2q3RYAo/AKbymty6IDUg3guPkG04DdvYmdSt1ss72UwTI/9cPgpT4r80
fvtMyyzANdDiAisp4iHaorncu9jddHz2sQymQht0oSEHjHFNCp7Aqn9j1wQxBj1VyLv26GSy2/9I
yl9RXpGplLRHTjVhCcjllgCCBLnRXrO9EQM8QE3aEJT2Xt+i0QD/yxxdgVVl/2TmZ0dF9iRivJTx
TfS8/hZOoRbwg0ZDV2YosIzrnpA2Oyzxmd00L6Gk0xQsc9tLA+z5rX7mL6J+guxszREsGIxM2XB9
99fZMOnyYZZigYi4nGSdgaMF4nKHt0pCc3WhUL7T0FJ4G06dhgidD3JKK8FNWbYKVxFohps/l51Y
u8uLB6cdusLv/lz7n9DPHWjfasQfJHvi9L8tRg3h8jKPUzlLR3nN0qAdFP+d1VHW3PFcEbzcA0vw
uK6VZogaiTw4l/eov7j/ScNtv1smqIyToan0kH89tqvKuYSj4DdOATwQxe6GXtEFxQnvFHAle1zD
vdUa+LH7INm1Hc5xw/6hbnuPwFAWsMcsA+1P47AI7JkpxBtFlC/T3o1o2xuPJuLKw04VCkPM+iX5
i6sZEg3bTdaiYmJqSwGwWHxd6vMVpSYeQF0hrXs3fRtwBRiENKKIsFV8EO+Bp+1Ov3/SByxfg+UF
m5UlXkDSYtb2k3nuZCUdle/qIjWPa/i+BnvuA+7oe7rola0G1MbI1F1K88x1PoDXImk8uaruvtjh
YORN4XK7FHSJXuFFmEwHYOb0Q6LXa3BLS+YE6uWymBX51Eby6xMgUBFLTlyidvthq23OzxUjulRY
ATRIAbiBHEJxdpTY4SF9ym97vpgZPjuYQgfKGtgcPaYYl8KhtqBoLR3y9QvRHV/5saL+/R93q92h
ZteYA44VYPsLvA2mYq6m2PfhB2QhuCmDp7FhXGS5njrbSPNJe0TWFRzCOZMLb16Dads8aLQJWCVv
aawVKkQ0vLVJVvo8LyIA0V7TM9KjuFLYC8szdJ2D5JSvIhYlYtwEIOKSDBAxocGEmWgj6l9YE3c3
4UiuaEq5cVZgZf+ytiuDzQDM5x1J0HsQE0cZz4uBSOggMuA288WaV16ofIKkn8suyvk+2p0eglLZ
6WukaNKyxiR+L83f5ik1Pj+XYbXCDpTY1etFQKYxsnbBlejpdlz+xl16OdmWYaYRGDa2exPysx6c
9gmqodZzxU1ir9NZE5iXH3mXg116r+QPHOKPNWDbunCce7N/apKcJYZvvEGU09odIXlgbWiyHyaK
tZq2BDg3iKPQYBfbzctwBpJO5CEvmtCWy3cxaEz9PhZNSWukDksH94NYtpfnTxBJMaknrb+NvFKP
j9TTi/gpQpFTMJ1KKvi1nf6/pLTq+CKTiFnzkJpIf+lgzQdSGX5Ps7QyfWwltrk8WKYcyixzrlXT
oXIpK82psnfFou6Uoy1o6Vg0+KePLbe+g4nlVuWvW9sMeb5rlH9xxQPaMxbl90lK5SK1atBaDfgC
vmNQvLiqP/4cUFXLiF7+xFafOUGWW7kKP37ilcJT6Qz4MP2ni9hqIfMVRU90rb2M27ZIJT6mm0qY
YRKYYy/kzMjJRO+Ywc2JEnKjY0D+Ruag2qQxIbHR8EPy+M+E/UK4++jSlYdtVC+nCs7zsrPVXhzn
SJEaOpwWXMd6qb5MrJIZajwjKYrphM+R/GPWCTA6AW9q9qKJtKS0gs0zzLbPY6Y92AUjDOf/aJ14
zOCf/Jf5ML7ATqJfQrdx2E+YN6D0ctvaEIXRHj0mDJXmrWGhxJ9dtcvfb4gS6UYxd1XHwyfSv8nJ
HrVsXi2GIUylgC53++Er2qD3D4Is6nkRobSmA7ZY6ZEcD/XDup4vXAfhq4x94UuQV0dwUOviUY0M
9opqHunfSzea+cv8t5P4+gm+xj16IgKpzJQ/85MteCnXFBSK+37hSY1xhrPum4Zx5LUDt5XksqoQ
zLTwMxuS2GyArDKDzKz0Au9gDAOJceX84mHW3ocph00JFYpq2fG+/b0kWqpp+RxTPGeepRcJln82
QdT4REMM64ESkhu4IBRqJSx15T4m1pZnI4bIfJapSNYt7FY/l7AP6o0xPVKqhfk+G2UPIQRagBpa
/6yeQCz4t2JmIGtJvHFOdD4eY/IRCFu0XWHhiRXKn9Y3zGfy5N7q78DaroxKbpWlNBkoJWsaq4QB
JwvcFOiMy+2uzh4Ces/aWnDQgh2046vU6AzrtZXxTSZGl4GNtXND1nR+wJO7o3Ww9V6jTlTJffb5
+U90l8IaFQ5N1fj+qd0TdjwZME64CdgUoLGoRZKXerUCX6gfr3pvpfZZ5afAeod3WK6ZvDGuBnbg
STLW+YVioe44ZRSUiQFSnoenqQ4zm8+HxHL6ceNHKkzALXcXp1UsxG+w3wm1Ygv++RkOfNBrQ8/g
gXpaHY4z3E+ljymZ67BBYlJs4rQt7p9x1yBlKpEb4zuIMWgQX4ii1wvdkLWhayQLm0iANWq3aIbA
0zAEPqH6/QjacBZJOC25lbMYjD7WzpnURSxOxxolYygy+IGi1diAZLdAUe0l8DpbpVOIUcLmTTNj
jlZ9MuwkSQyH5KZqMFR40Ho2apKGspKXahAUzZP72O451bMN66yJBuJxxyBJM8yiT/0GQMGe4w+O
OwVKPiDWHC3BRGr9QB/XOmqfZXFpM0DGXN9xqj1JhiWkmyaY5lkvh+G8G2Q23ua5rBBO4yYKdu+H
ob9DT/k3XzVE5ETGpC16G3EKUHerxISVmDBFk8VkLRs/wxocWumC1ot9PdVheoy9dtkyx7X+KsBP
HaXvjubtUTpnAVZCzq7wasbxDdW2ZZdbn/TJkh/1T/Qkf1ziqAm9hOV6dVy9qhmKbw2oaGoXTCLE
zJ4LXO8b32ktezngt1QkLB1nGkyjNTk9lOgeEEq9AbAOIgcgJrn/a1CMBMmc8xT+moD7z1x/Ru89
NqjnRlwtZIw9HDrELCRwruCvwg6R/bWEgW0g8I4b+A5YDvILYslKHlXEakM7bEzvj2oVnCs4/zTM
msBZQXLRJZGhPQYt5bdDbmY21PmDdJYVZlfX3VJ0nC+VKDgeqnRVTRI+j71dQMdye8lJCwSaF+iT
dX5r22UqbYYvPW7RAYbK5yE6a4l010Bj3qCS6+yTP847czOGB/Y6vAgpp9Wf8se8GuTdkoPxHz2j
7A5XW/VdUn3EeU2jNmvyg3+/MqtV3S802G3WcV8e8nn7KLFSB9k3UjlBa77CjsZAfJ4KnHeDMNf3
2xVjPM4ya4POaObrfRw/d/AxVi1mJLrmq3Zk6ibsHUjdwK493nD3wfy4pY/hQLXJS5OolcTsbuZF
gWj50m77kNQO1xZSOq1OnP2rav9uHwbzZzc2o5ljD7rRcfP0qN3QdVA7UajznCEVLynGg0YotHpW
uxAoaCpVx5WAiQWjF+gyInWsVu/isaO8d/JlWGwo7/Xnl4x+4H95xODMvQDGvxWGIjINlS8+9Gxz
3jK7Qddj1KDS8z1XIdPMlypPKSEvbaqotcxQho2ZNAz8KVZzxhCecVQobh58lNmkplhpAIRW1mPz
3SvMEdxiOMwwgmuRmXbkrdZ1MZfqEEN59BiDrJ1RaMgTJlhQFVjHkEMg4HhfkSbRxx8+FH7e/Myt
PKI5m32PKJoISBTFsQHEk4hVESF09XAsQ1eKj7K9aDNL5IJQvVXqUXhDfp43IhNx0Nq1lBgH7pqF
4S/zZDL+RF+KHYh4ywBVb1oEebLLwwmpSRH9c9kE98tUhtRQr4UZVxFYARNbNHcjE4tHsEKo7pWn
aIcKMXgixZgRUdjmMJmXzIpsjz8PJB47uS9TlhQ3jsj+RpJlQniCVpfAGonKQNgrvGDNo5nJqMCM
Jt+pvuh8WZD4660k8EuVcAUGRf9Sv+2lNxPYdgvgID20lQseoSkmkVSO+lLz2frcF6UiOyAfhcHj
We5aaJg3zO4nbtQNzelLOJawdOlwpRrxVEVB2D4a0UtyYgMzt1eUofuE8cmjIlBc//TDIeaypi+2
0291zlAxj0anX+jgS0U9DzYqRWVs7eo/N9wP8R5F/M75NFs5P0PEmGW02MimCs6df65gOyZM46fb
qVc+3TFbUDB2gf/svqliS4rjvJCtRPi8+F3ePyuL5XMz8JkeSj9WI1CB1mqnSjmit12q/giDN5kZ
Ei+OqEFqU9LP+yGkOo1qR5TcB44yOWoZT5F22fMm3kVqv48XwqSPWGY4yyTHorlfo5CmmtQNepq1
Qm83Hzkmss5T9W9NBkp6jBfY41rdi0Y6/Mf9du1WhJMmBXnNDW16HBIFAmDh8S/P/hxMkd2vSvp4
AfmusbnM4yCb6/NjRWm8/HIvMAB7iPxGVp5U4Rw9sxP5iFYQRcIEW4YpTPo8xFd1D3pOyUe9WRXt
1Pqf3KpuJnCnpkFLw0+65EgQbOIZO9fGI0D8fYVfuCH1WolUCf6BbQd+UX2Lq43eXHxaPnyNc3SI
HfVWiGH/mH+o+gtTM5aGwdEDI6x3OaRxnQ0bU7znxbTf/CLBE3pWI+jcRvh1fy49WVhK4MdDKWWl
IhUeCjqVynC2YlxmIAL7XXvpTQ16l13zWzQgDlDnzdNHfjeWt/1tHUmvJWGTHmaAIjTh/zCJP2dL
Qk9iN9CED57MeUDat2IAPAOsQcnUaF4LTZzfUvpRgQFW4zP73QDV7CfhUnv9MRS6HPabufb1/tY6
uu+GWdcgIkMGEXwrItkmDmQU9Tseh0M0nlUIojJYIe63xvNdB5KIKwGL0NumnOH18K8ztOwiiC9Z
C+FN8td4kfMKewzSc4uZCEn5p91LTVvUOBJLWl/7JpIFiVVZXW+qRd3h0/upr3TaAdjbKSYz+us8
EJ+8DilWyiSmU0sORMaW/e83RQK+vQ19mCjR/2tgZfHK2cCYw3694yHa0EvsjfjLrwrvl7XwkBZn
i6RPS2jp697QkJRo1H8sjU6AI3aVqiUHmMBRYCcW7YOXnYywBtFfyOAw7BueiOvMC6W3kky7GgMG
cTFhzjmqheOhbGnem+Z+dmp/wD+NpPQuxnCQyjkhK1HPQ2JysIrUL2sNBTV5SF1NsqcyMcEhjhGL
kgAaEohM10PPwdBY5cFDVonmZ1Q2smgIurRQJ99v+VmIn8BsstfRBTLqwg/sUzRtRXlMit3aT01E
0yy8j5R7aUAnlOh9//jOcsv/zIIQT0D4U9ARizVlChq9/EpiMvc2UHhOli98sf51e0nkNUOZ0M63
mOvCrUvlCRZh1KkDkGqIHw6+Wmg7ACZLsTy4GwRZWRjYKgijxLLNc+VZ1pHxC4lO+P5OSzN4FJjp
rnscMMh7sMypMJDrtOYB3vZwGT0HSNtao6pCaczKKOwpIoVZX/XnlmjCJYgOmfCX53MYjmfT53HA
wUFSIrDQmd7LRTMsa1lnnbzB+zPEldWWkoFrWCkVzFcYw7wV1jgMCnuIFGDOw/8BESs8OqiXfkvF
DY+/4luEEIHxeVF3OEcMlzfDEafChlcwENbZpMB4i1YBa0VdmFOFTUAJeD6zwgZSF7D4u+UJX6Ek
X9KO92yUWTsqcuFQ1RVZRyCR+R1L5NSwt1m+3en2FiIHiJmPLMPExjgTpBBDfcdojT+psgtXr2jw
usv1r3tls8WYnL3/WcCotLnbQzrd9la1zorUERljSxSsOOTPr3C59/Lxp8CE297PdX57BGs6WWrj
DC4+Xbg/1BVKTyIFVB+5onLpn5noMFiFTZ+ab0BbjiUDCCBCP0MKxFVFaYTrgeFH2EQv3++b2Clc
2XgRmq/ZCZSaYd7kJAyoGOC+kAyBTN5hMMLkniUpbVRcfPcjsFn43fuJ1bHH/M9sO+z9eui1HIVp
lZTeYWfMfEaeF5WiMoj1a7zNejTv+RPc+g+gDIrHN+vNZIXVnYCREO57c++u7HWkogVBaFt9OeZQ
qyPlfbsvFRrTcU9aLDo5+Xd+NHtFE0GPi5ZNP70NxU31++ZrtsgefHT2TTkU2hGrSeEmAJtGZjFX
Ervv5hPykQT+rxthshXTdDCu41+VhEMvr9qfbEZQS5cnZEMQ+646eOT6TQ8gVllm5tSDnY7ku6rr
/TjZs0/OsruBS1nd4n/b7yHdM586GX4xlIO2bNWPOpAmhv8DtXqYO+I6RPBZvZI2xPwwqa24mQWJ
LlmTH4k6kI+/WIQK5var25PDogN9IMm9UBkSsTSX0GBW8MvoiClQ7r99+ZDFO7lRqWj8DVUBjsYP
tvE/kqoFc0ugOJq9zXb6sOxEOev8RMXTeZGkI3WbE/RugIbby14nMqM2fosGXYa3cI/QChPEyihW
mKxUIyc1GGy61S+Srp4qbZPVam1kdh51fs2wU7/q8zIlGvtPZVDJOe44a6kdihjVgrI++79CqO+o
yU9i3crARiFvCALN7+CHG9Fg1WKdrYdP4C8ISUjBoqQ3mmeZQfrGo9QRUQcIJ57Pk5SbXh/Ih7gX
6KfvXzwI2Z7ZSxP1+o546cqKUBxL4KmDpzlO0rsJwvA8KQ4/gmW8iZbDPC/cvhW7SmrPyXLZ/AQG
0ocNkWhy+D8Dyie89VYoVf0K3BFx0T26dYXw7tMMxQjAb/jJuZN2D/4C0Bjd85zwSoIMIY6Qdun6
IcC7BU68gSz6SgEohUmniNFx/2lEsOEqx++aQp8rF/cTY9coj+N0nqHDS9P0LCGZmb3Ax6z6wahO
0nnpurhhyMrWuMnNm5PJHWbHf2g78oN+yVZkg1cptEaFHElaTiIkDLJJu5fVO/P5TeqWAs3uzAoB
zUbPFSQtKCtv3CbXKBdyc6zu403Tj3nMAgUdqOERzW+t4z8T0WTmVmnKQex7OTMOWcDAAXrr/5xL
vaet29kx7feet9rwT1oNKc5Daz7hev0+vAdVH73KTGqfDFVIzQrLsyGH3YaB6wKPG32X2/rxruqf
hWOjGx8DLrfR7iN1/BEAu07DBYOP+t7uBB7hY3y4nTe2HL49L1Dm4dGI8gcuPtfEtKe1sl9iHlQl
Y9dVTKsLqELgNxCCBc8V6PQvw53uoPUlt/LQQlabSt64YZkeIpRfWk5ftVmEMKKjfFyAxQIQSOE3
finfRs7hhSvYqtNwHGO7C0/XqT8aqy8CxOSd/muV8TBSN/F/4F5cl/k6FYJnj/sPZbsqJ3aEvEhl
MiA8NjlWwefIq0agdBTEYDjYRSgBm51tymdHu5Z7nX9PKn146bnR260N9JhMJ8AefrNx7peEKfRn
Hfn367jIYgUsUjaqTVCpZQ3PM9ELkNmepb2ybAOvzYCTRXESk26Gae5DQNjCA9b+5X3kRph+Xnor
koXF2BqVHYztkCtL31LmLr5vGjLczPckdwN5sA/4y/ra9iQVqnxRjMNKXWmM0fMRbSWC+HOwTUth
KIY1pCY3NY5rBXjhJKyMb+g/SXMQRnyWE3tdVEJ4C5MK0E3rtNl+FdTj2ZE0TN9lZm3a0shJOTX8
W4CkW3Nu+rPfO+h7j8uBkYOB4adSQmQP6narEVIYAL4cWUBW89YzTcv8uk8Eb22UXPDd4Y6BdlRb
kHoD0Z1b8yyELdqs3qBs+bgSsEIwNwbiIf4B+PWZO8bTXZ9qffz197AXc4jvF1egJSMARt82h4yH
bfZPuZeZLH8NPy0RES/en+StLeg4ZUgJrVu5My1JOqnB+WgFyhlHDHrEa3JNSjX2GOkpSv+B4aoF
TLqmT2AFCQaQnLTHMrWGBMTz+ghwjdZdoKGOnj/M6xgh7P1DGazsHWsg8JT0ySRTYKvJgjN0BTT+
gc7Ey+e92a9miaRM7LNi4fGvheTBRuhNGyHmAp2sl1yvvvpXZNghkH0FtRVghRNhuJC5qpApI8k5
kzlS/9LTJ0JKKytRCgju/3Gq3AsLZQTVbjw+543b9fYWThI3cbj56rfQ+0hk2vygT6C7cirquP/N
o6nV5T/TEIvFE3B6xoCXLFni8vkEhl9/q1Npp05V0agh+YU2OR88zF/lIJHkN9x7PLX1qUP4KnM6
gqRSsHT6ZKvnT/A0sAyDBOXUm/FlBmb6MJg64IHDMHbtj9XKFHS4hQUKUnSVpqIrf6jDES+V1Sm4
LSgQhzt7YIZhSgDp2x/u+gpaDVquierjdsyAiUWZDkNS617LsORECkEGjETbBSCPMQlOWoa1Wfi+
yVc0Hn6hD+BTFRR1+iCOwHX6fGJfS+K/4fcVOs5htPN0xqt5G+UvFGuTRJBoqiF3KRiSxGIBqhhU
Zb+QP5QQuEN3sRXkFY9+6MIX5FoP7jr2j1YLd4FyEW+kp1j+Lm9jFJHe6l33lPw5eUzOrg4G/ZHs
8UhW4ZL2VbWyUvJ226yS2FOF3HD8TfZcoEIIPp5KlEWD1dDswyViT/vk0FR7vC42yr8Su42XPx9K
u6dHIh1IhrgDHkL1JRuwV/QmGr4MITOjOe2/NFcw93gbgw+NLZyDzrHncc7R59CWXSEaQli1ft+u
UCH2WbFeUP22SEtUV31sAkuM5QQ5HSGJyuJf18KF2UE5iEOJR+9A+zmgcDCB2k4hQROEjsOIy0HK
u3iLI/AFuol1cVCLxIdidtV6V/s3xFqGg/C2RVNF0twuMwiC7qAs33dkl4lli3RBse++czm9TKEz
ZD3aozJdoxAnG+Z71LovnCW/dsN9H31kBAftFMd6kxAbaEz/er8P4vVeOfIA4IS1mwA04pMAAaa9
UzQFTO2CxqTXDVD0a83SeE3JPpLgqqPUD6YyonqUyOt70CpVfeBWcJJNrpOzsNYKvBVXn1IeJ4Mr
++s2DhIOXkw6fop+9Ffr9vIpJQjQm5Fq7aWxAp8w0bC2j/1KVTNBql59KMY8Xv/D4uJZ7iFX2RUN
hN+HkCK0UCpYWsc5ZT3vybH2Ep+zpH6rkOjorOsEM6JFDefscF+sqRelawGMc5Z08mULSne6safy
m3U49cG0Iwq6FmVpJ1OkejL5SwE0BBqbOORpY5cKVeJd8z8mYUwVBNt+MUkHePWR5ekLN0xqJCUs
BLA1BqTXq3py/m/I6GqPGtFOCaQp2X3SrrhFK22j6u+LYgiTvfOa8budzms4HgdzIvT5ZCTeyIZG
5w07QkdB8OpwQpSWzBio5mfEg3gpCAP90/04lO8u3vFRANmmf/zBv0YF/QutTn5cHJ6Y3FKhPtu5
M7QhBgffNOGDgg7AWV6Ej2Q8jPrzWPSnk7dwtIfZFm8hk9TXMA4+4J+EkuE7aKPLAdS9OYYDkCgk
1M6rehH5oU/NRpU26nCYiFRMLa1yzbZsLWnsEse7x7KOzEjqaaDwObV9xqLQ+Y8CFRWboe2OwBX1
UCz1IrBkjBgHkg2tm5wmmNM5tKj7ROFvhVPwlUFeXbgSwpRWF4hd6HrYy9s/+t6F3kPqHmXzYHy7
Q0jhR62cQdu6uP14c+7oHpzWY8r/OeOMq4mcOYr705ZSrhmD78IGG8CNAlA7hkyBNXUlZ3jhWDpW
dcBrtEDs/ViL0nH8Xe1Q8ESY+kCNwlWLOU2BKtPsMiE8pIvLch5cs9uYOOG1LTYuoYB8U+MjL/6f
2Keqq0Nt6+5OynxLnAZEJacn4EcTnMvtu8gO8pecDjZD8Gzw4SDYXW6fO7jpsxyAmst/bHWJAbVh
u19NIFHLGQd7f6G3JcswZ9nnzW/75Wnbjr1R28i/0UXokdWoXT5EplO3q4wyEYmIjE8cGt9D60u2
R8MGboY/zqsFqYPEillj6XtUZciEWLln9h3Rps/xlO9fc7K+yny03Wd7C8X/TrAr7MYlZrcYfFwj
RSOaDID0ZEn5Sjk7ccjLJrkKy5M+zWzXW5bBLW4PgH6N7nN7fGm5xP34okxvo4Mftk++2ai6n2Iw
dBJUhiTW4uWCMNrF2ZzDF+U62n23Nm/ENRfgW6RXHd5latC7i/BjCLTAUBlvilLUUZGY+Wp+Gqus
iGDfCf39uoJ8mMGymY80xPlXZc4HwfnilhUQkyPjRK2LIJx+GDaDdamCbNm7Wrsq2cnIr44tFL29
b/s260bhGGxDl2dSNZ2jOtkuh62VR0SjyyKsGHNVkQKYvRyhACzKEspI4b7nY7mm7u8tVjEkPR+7
EU9hCxOQNAFL0MWvNTY/Pg2mDPIE8ymU5nUy391tizpxpS/2RzL1eIQ/Nh+EWYAwgGk/NhtI9OQq
yPI+vJdV/+AIAjz9n/COCP1Wmse7kqGAADuHL4MSHYEkGtdovV/rOCc3ultNBh20QAI8xlqRGuzc
qpvHniSh7NRcDVffAzlADn6+ixsxZpx/4/vv7SwUWJDV0mlmGoOnhCEHLPgQV+tNihbKEgHTeJi6
tx5rUE/nY25lFsVgopVohwNtqWGTcm2NqkvTlQjlDkAUr8dJtgOJ7eFRxKzIm1kdMvtnWqkRLZ6w
FxIR6OKbj5LL+T7GgLBIr0Lk61ai+F1Rtf2efgdMz9iwvkZYe5lG8Xb6GkrE0ViZEJfjY71W1Qzk
xgZkWrA2vXIwm+gFgZfJUrr6V4/LPTzfnGSpPjy9zM6WSyw73NqgB5xzBz4YidnOoUM6VEvTsqfi
rhX0lJ85Nbe89UIYGJ7sMu1svmoNzlN+KLCXg9LtaLKs2lt7dItp5Be/JFrH/9APEc5wkOr+Ooe3
0IV/1CcNvTEgYWy5A5PtWfKt99gLxhpiR1rptMdcCfw+11BO1mSCTAC3QPmoGozdCaHY5u3k8LCg
MF+vr2tc/aBJ3HTFGx7NtkQiRXYZIUMuTneOQfuC0XljWhWyMFp80DRc0oDnV4DTCWZHiUyEIF56
kZbjrQCuhoHvKAVXNwW7FQtke8rHSjT33tM4BI2OsA9P0PW5NSU5IVHttg1YNb2MCkfKSg79pq7n
dfCPpVdjZBuano8CnM5dAGZG0THfR/307SjLfEl+eN2a8o8EwCZL+aIYjz8gXtszNXmipzKNLONI
QFYOgWBKPqF/4iDDsiocFlpIXcrOHRcap7BQWqTLz/ufQJ1OC66ZQPTMlQ4MVD2BNN3gWITEUDiB
vmEODU5WuCR43zpXVSg2kQGl4VrLweqwoApb+BT2PcI1zJ7K4lcdZqijHDKL/MKLxwP3I5QBOb9k
7iiJCSBLZiRMG1+/UF5W6/hQugYw7dN+5fJ2UBhkuA04luC3KM5KS23DEMur1HlhXPwTIpdAtmFl
YBlm64esJv52SqiALL5YdLEmyWmGJUEYeAHX3V1vjQhWa02DfpnsueuD4eIKotA0a43ytEwIfSPi
9MLaacFmwdKr0AbFzNavT0XlCCtON/xlpt6gftWAM5t8ZUFmD6FgqnBkUK1eWl0r9O3jPD9oDknR
shy2Rn1IqhZ0c8H076FpY1RuhMkRD0UeXI1MHNMcrAQ/IyQNBUTkl/NSUgirmT9PCdzZHmuDME25
6MY0XhhvgGdxth74szJCrxvbi1nubjO4xAPbxOqaNz3UNQMO3VCnnCOJovOZ9DACSgNYdY1Ae6I9
KxAjP1ERyK+GJWEbp8WANJLHE7H2gVWP28qJADGnB3mJyCYKTCAexwHlRo5wmAOg4q0oPjKiBYJH
zirLjdImb5CtqvFJrasMwtM/752iyUGgULN8or6Q4ZF8PkNx5qK1KrEvvXUW9QMbjD4g+xDq9QPj
CH9LT5e1LFBtdsFJYt7WveqQeWX2+hI7W/r0MNy9wTcm/cnzKI02FoxfT2dK99UC/Ob3DR09vdSj
PKruxYYS5kAg3xReFM7NRHoo54XqEca6366Hu9zU2HU1pvdYBFY6EOWh6+aBp0ftY4SSbEf2OwgF
SwOcdXbYgtuHE5jCcRQRLzgDEu35F5LSgxLFSxW7QsIuZjx1f4EZS1b8hPHwLzh29dlPW+Q01tbZ
LJP3EtGMRtgrqMku4VAXmPVrfvPwa4hV26+gGoSSUGY+vRRIa/kf8fw4KM98nkVXzrXAMApfgvgO
L5rI2iaqnIlNtiM/mlD3WNnUehdq9sdIPFjM69otfj9dZkC/eYDY9QZ+52I45MABPuAifWuzQQZn
VIwKJjdwl7t6V3z+IeGNgYnGXgedG+YYf+4K+iRvwPLdPdAg0oFVJYAnT+bSXCBPvTnmUXTRBK9s
zk1dfPXwrKlo05AIchDUSZaLl0tZZeV7nkh+/VbDXNnmnXE58YHUqiBzEM1qDNQsfnafz6Os+8UM
vzOS0eOH4bfP+/seRU/JoxLqwsq/mGoNBHyi9z40Y1YJOJ5iKCFs8IHEqIVGoO3sypff5ALt/2eD
nQVILUXI1uTa0ywEbAPnyYUi/VeuCdj0FqqyuzzJRVDJ5lkF3fh8VLlHxH4fMtPk/NVyK0sFUWNA
kQ1BqPAAivoSOd4tAMwBbozYCi3WQylnP8tADRyhUOC2ckREk+GHXYDlLa98sJ5xa9azYpWCkDRr
PoYay1haNW5XDySe4Cg45spkOguzXIPWiurmh5+g4kB5Dszit3m6v2cKMaV9phC67+DORmxXzW2g
5+pJE1KYBnaxt9n4b2n7W/HgK9/8wolu8UWFIrJnMfPk59xnW6vGhNWEJN54KdlD5elt6floymRo
C7gv1ky57+ji24WJ/1hFLM72BzdZF/QWY4M0M4tgDMui6Z/XSvkcsKLrhhlcO5p7Io9MIlsqJ2Nf
RJIpZPi/Oa/fc40gf82UlCTTRP0vU/bUABywu12sX4evauqY0nRj9Uw/md6IZXlSneRNywogQD3e
13ZtFtm7SHXuS6lLEEHSN2+PuLTXpghhzL/5Q2VnN1/cZ4peBFlMOyzPjzVGbrz6CqA97AMTrNAT
ZFM4Lmn7iojFkyLZDnwCRR8EKqNDxjzvwmzqU4k8X+XZw3PFERGLf1RiSawnt6Kz9AHl7fu087pT
KFeiqaSa5UH+z4wTWovcFYx00aJEsOizYaxrT2mPBww3yHHV3tnRVn85TKp21eumFW2MYz7XH8Ae
v94JSbA7SUhj2hA2BaazOhva5wgtl5CTfYnGzOH14YrO4IU/hMmIz1QBqiBOj4/ffgwzTyi7B41P
fHHpGbwIe63yuHNsTHpaQ0ODiOnL3X9bX18CLqETJgpHbTRzfqcC8qqvAPoCCEBMGrV4BMuDhyJu
hGnt29/Mix+42CxbNE7PelzobzWcK1BJSfPOIeKVuLb+frr/xEnqx+S+vs4toC1YPkJNw5/dv+Qe
6+K400fLFBUa1EIm5WEjcGUHTt5V1RazJYyef2NMK+DUq/VxbYvPylQFBmWcchpYydY8rcfKnNDc
0hV8pinkxqppLPeyZYjMLpfumNt4MmZgMhDs8VO0qt3w31gq1FZXNCLjtwXEYj59AdhlJFxZNKEs
V8ci1ykarcTg3GdHvme2XmNhEi6bc9lbG1ImdOZshHP5EWw+HqoKPu/cYcuPOcQNHjFN2fns4dRM
VaRZbguBIVXCrUoXeBakJH7Kr8GOHjzfIbCwLh2dUzvPJz1szdjapY6cIYJIk+pNruNBzFdwon+z
8ObImQyIRCX7kg/A5lHecYDWYjbdYOlyyUaXei2Tb1ezLnl4lPfeFbWHANz538NgDAM9hrVtD5dY
NcDTWMxblUubSH/qvW9TmpdYPathQCPj82D24aiucmUPGbR7PzmBqSjvBQ40bBBv9LDxPF9Nn3pt
mJsJGf5L4o1KE2vkyhofJkQLjeGWyFES1dgkozx1ScAnY4+xqAoUHlBjfO7wz4OgZDtqFTYyQT4n
Xtk+U0zQ8C6PTqO+IHWHfy/Hbu3ZDiixdgSqID73hOkmbQoLUZ+N4f2AqXNiT09a6i72TZaQURJk
OTnNSSfY5/9ma/AxFdIEUOrPcmudWDPzwn+dR/K6HbGYSIUZZBbhjlMfKxJfRKEqijcrQPr6EiGv
WZwxse5SVkAWa0dTijaDPGuz0f98U316lNwQmr725XZrvUM+urh+U5yqUTyeLEogSpdBHpjwkWYL
nI62oxh5vp5GTMOroRJhvImPai4GZ4ZRMcIsZQOlk5nTIttDwgVj30kayrrfgaOgPmdJSqg8vMUg
LgTQlY6etZeE1zeI8gLUb0zZa9WiWSEjh2BS3gEqOkh8S69clw/XwS1ydLx8aIl+xI2TQBxcbmKv
RKqZ2tQHpCwfLwGGaGRI1jgf9UMyov3JnGYYwjLwc6vIg57WxHM/vLGH1OJWVNpYrgs1wI1J5ElY
kIBtBKDuGG3RXZRFBRhMJpvbl3eyE1t1ZQjwcAy+m0zTtUB4bXbmDXoJHFFbBNReCp+eTjj24QEi
ratJtdNcbtrQ2g5MtV7YZY1vRd55Shy9q17l23ZGWUqvy9tPULvXkI1cgTTXvIUKX9Qvk5gQRNil
yD1m9RuzdblVPoubAbKKIqH+OuvwYaCzjT4K3XWXOXdctV17mSjI9lHkaM6FLLc1H3GUdut2n5E1
W/j0LcbdkCkeedfrbVoiSv0dJZWEpxuL4BsM1CiESCpKDf/Mkmb+zItFnF2/UK0NeVvfsje7xzTS
9zhBQZMZmaLZrVw7A7EST3vZdWbXmjO5dGFR5oT2rz8mrOfSmXoOSAD12HSRnA87G5WJJaXuOrgo
Mp/Srj/eyc51v3+fNGKXQEDOYq3AYhEJGt26wmNR2U+E4fbxc98CkS8xbnYorY4AlJdVPQQaE+h9
sz+BFHgEOrUYqLW12ETUubSnsjjtn4UEn974chXLLokd1I/545GHIQ+DYS6Nq4h2A6GlzdqUsaQR
x9032ZF5g72Jo3sldILPR5rnGcXu9nQjIThjUqAC0aWx8UsZwLdXOVsJ8DwUteyWImw03F0RdpQC
51PjSnzukfJ3zDXdgHt/xZrxehSAc4HVlstJ5/hFmz4C/9MP0gcLoq1UzaUG0KeDBdrBUq99MXHr
Q0Qfc4dP69nBcllbentDfCV96bxFIZ2PuBj0wZ4MiXCTLf3wiFddpJuNmgD0v889R8rmDBkkfWNF
AK1aclQ7j12rLxIaJUd6muLTPOAOfB1HP9VglPDvtxY/GtNkazmVWO8loOh+tvTEGbpQeqbDT0X2
eqpZJguv/9Z5ld2HPh1x/6yPIXs7ALYnfTwHH3KiouXVjv177A3KFfV/76R9McbQTjj2mlC789EB
10i0pNHFChLaReLavGeODFAod+5G2He55AZGOMdyxy4JitxA3ofEgY6p5wtCBWBOjr6led6qGWsG
9YP0+tTBOH3FkdhvQ7VTMOkWXv7083d7sXeSP6gXYOwpYnkcYp533WVuGHXCbaFKW4lWI14GH2Ik
I1FnPt8vc7bQeo8vrJp7SL/djCGY03XUDC7Vrw+X7LES0drEfJASXuvX5Rb/q1A3/gXH6lVQVE9t
v9NCYVnq7OI1TkUeI/jIhmaSgfcA9H47R3GXcp/8RZzBvPo3EniRo40z8/XT11ASlDvK0Ey9vCoo
MU5xvnMUMc4ibL17SB+NCReeYbm/YszYwQ4Q5hVFDM7aE0b1s5eIG1V1gA/Rj8JETQ0D/KRZcYef
OiFC1jGMGuiqPEsom0AwG8QZkwDuu0wLqMWf+psVmigtcy0rhfc06B6zJl1nUw3CjLETKE3hNI9S
fEGacF3B2GBJSPD1am/qeyKaLESmyNgxKW7ivpLq1pHCFRo27UrI4oaLZJQspfprk0LJnONrXKo5
EsIlUp10HNbHUantfJGo16KYCj1nKLL1O+h2mTTs+spBUYh8WGJExOH5jOkqNGi+80lU7z6b8L6+
sUGWL8XD4WGIazcp6d4Pew+/jDRHs20NjYj9VeMyIbSXC+cnN7nmtc25VMDBqbvu429zrFaOCnCt
6gcXHhRgc/yiGsBbJgA+63O7yTZ6geqExfoauqgGawwOip0mOvf+kwiTOyKhBYZyjH8PelZEm6JT
iQf3zT1NCac7fKqLUDzd/QMx66biJVeIDC+KJr/tkhlkX5EKPSWLAWpIGQOq2JYKx2r1bRifUmXQ
6OBSe2oHn9g8iA87mlpI1coCsTvCpDUizt5odjmpCTO2d+NbBbGkVPofvDZRPV7heVpGjaP5nnUq
5tGNpGVV3wSNDYigAczMAyBLmARxROmiPv7w6smQuaeVd8EkunUSRv9f0X3sXGVqXcCeZLtd9ZbA
WaHLtmD+5deSdKCvOouSN+EJzUFeVs5TgdQn6cHVjyhXAuNMfnAir84bvbd1Xj7UgjvfE9bYGLPQ
V68blfHzAR9oiffY8HP/7JmX5eWhDwo0iqVzysOgTsJWQH7Q+kX3FuESl04gSyEcZA075oopnLgu
dPBF7EBtC4JvSHBW7EJ4U+WFItSWlrWsXEeI663lDpDcgIhBM6Xfr+MVuHURfWFwbeQSQzVuDNff
atEgvlbkOfOSLYE4yg3E2uRejXORN02cSmyq/4Avdx0XXQFhRQd1yKUXqVbPMAzwKwEumkYzb7Tg
NpOw409OZrKhXTk3Ve+AdY6w5P5EE/pGskeqidZ98Jx0ZbsxQe9WMER2//cy093lzmec8z1RO6ar
y79GxuuWJe7kaqlE018PwSLeLFPzAqubeDSXBZ9WKLKyjmUZnjmCKbJHYofUzW6ws7CXFFn3dq4n
lwd4fXSLpdV8Oh8ivW1lTjeYCeeRC/MxFXnozvGC8Gx0ncSyIqqAdUBId7SRbmfQQyA6RCFxs27y
6fvUJvovTDhjTsIZctaimiB42hRwSdZG9rH+UbRGXhZeHgv1SSPYe9oJS2POe47JIYXKrUeWTnHw
1n3zy/tL0RfszZx2ORNHlLoY60HX4iAZppZdiPdPB8tWKRZyy7LBJOdvEJh27O4WR8rImE2HyS+l
/SgQlx8GRfsxahwTVsBO3mIJt1hg8nx+KJZ040PyimQZq4qTUCBFTt2+D9SQzX6tbdQzkfbDUg+M
aRLkuPrwfvu1ArYQNy5rdMTQCY/2RuezM0ohmrCwEZrrZ2b+JXnTpdySOPXafEQAnurpI3OZ7isn
eFV1KDSm58rElbZCy+JMuepXU6dsngMsVwHnYQwTx3t3FLr9VIv6qTtv/Pp4gJ5wGKyXfj8eq2PS
vemlTqTnqmMcBNFDFIIjbzr4LpEqlE6s2Ak4Uw1QNZEBCal71r1r4iCH+lXhWThax8CQ5cNCw8S4
opyuSzguJcr2gTw2WhnmsgMt2YXREHGOEimxd5gykm62kcAVhwrHAuaXI7ZOHz3nYQR5MnQlrVqI
Kc3kOPPnYWmTVKFt8UH9qJrhXa5AQpnLpplM0POOdBedT0Fbtv1sY7yFpS7A/cvG9oRb5ti8PvrE
FfGEwCFk7dmO8HWdq2UavJdPIQwIW7lt9VeWsTdMjwY1hmaerZUUyaDE9+SzeqlBeu3nrVu4zlwY
4VKi/a2YRXAOIVn6lQjPGnldc4L4hfFuMIXaiWXXiI81IOXne4v2kBEiDCXpZlJBjuvV04ukq5Ms
4KOAxJ/Qnd/Hoqawv4V0is2+qORSja4lvMSE69fVoeiFlcbeCHXpMSoOId0jY/lGW1PCZCm4wk7L
aSNx2IBBbSICHmdEQwPCY5+FWChsHgd/9CpFeouCLbmBlX0SAojxoufexNGeg4sjZeVU0gmrowGH
efmu+AIwxy05wt0RlZA+o0cAo6AK3iGylHOuCQxwGPEhGBWiP44nJvkFNc04nC9Ol7/VkSujHJnt
UEGgXUm7wS/he06oCuZ57W2qLyuYK17iBcaKR2U5t4pBuJTIn+qwgRCOtW/GH2v/eCAEkIgAVi9U
0DOMMCzllOr2nWRHe6wPMFZ7TbAzzRQrQLEWJSV0Dn1hNwJo9SR3o6ctsIcBl1GhTStDuUHs+p65
LvI/0grK5jeYGP66ZqOwjGUvAbKWLCliOC5PfsQghtP3Z7uaBEEUraQGjFC+z8v+8l0OHrtX/hDa
ASIklAw4gVo0GFIzkLlGiF/Hy7Ki6X8lF9llVitD0qCcOuPwWk/I3P6cOBJy/vrek8AJL4lMqYRo
l+84agWTYzR0k9UgbFxrFOaOyO3b9gxvZrjYLv2cCYaAFFm2qXwWGBlGaIzLfqAFtc2LrKE9UC9e
SDagx1E/O+6OK7i8qKBqaHQIyi5O3uHKgqmqfjh+PMQnIgVAyV/5ak9Q0/PIGuqjpnS+7cS94+Ps
/ocm3Zi+BccekFypd+f64DCIplAVq/VAsKa3y+PRut4OFGAuPg69ANWXh31FGbEvwPhcy7cbcD1y
486Azwsx37cFtilMZnW4dGPgb94Q7qfWetoAi/eBNwC5OkHEUyIILDBLh+Mk6xriE5QlnWiv3Otf
gwMBbtclNTPZ/+nd0jJZ2euossO9Gu0QGzPbVyYZsSCV4jstLp1/es94i2Xxzjt17N6Q83wAtq1F
nnGR7mSv7Jepmy4EqBwyLYgfzMsivuui85SIsftcWZs1aIR52LdK+p3NlWY3dg3iDgUPYRsBkJg3
ZWEFV/PHFqym56QLySCPf11qHjrZS7SLaTvdbiO5DmhvhmDFnTx5PqkkI6+xinSZq+SH1x/VRSrx
J/5gCoS1EpI5ZZcYtnt/3t1ngU49wsQDMT0neQtf1N6FUODMleRkOmkFcXkjN8ZzSJNlpe7gHrqH
ZUNl1Ty7nj46xiSGxhAuLuOMiV/La86WIaqjh+n+CXDAso5xgvdmOFysDkCsv20I/JR7LMaaC7S2
5a5ZUU3hdmfS7vWBYCAjDJz01b5uokFDvkV9RWtuno+CaHDRfbrn7A7I0ktYVG1DttOxWXE9oWkw
wX8kjUn3wBhgzO5qNjByaXzo/xIdJJ3K0671GYtMrxVtxsPQdaQiK0t8NRRCmaHOrxruM9S4Z35Y
aq1kl8ISaTRagySoonXAMk/WDmi+ur1fGz9hphAHUZph31BqjskbeAQCq5r195sdjquyRpKjUceV
YLHmGQruicHkxWwj1YVEYd173WopUeMtb6rC3Rhhgba1HkKvm2AyyWWYby9NV9vLXSIkY0rWTZGO
iUPUff3IvOXASjIMIRZUv7HYzSfeM14LKCzmLw9Ez7jgqqzmvjEOWYSDcTvuEHFuA9FLjtlMUHsD
UFFFoua0k9sEYg4ISN3fZH5K4cE6+EuQdadII7HIu14U2JJo0vvcHeeuquvVkSfVJDDwxke3u5Cn
dQQA2Mjn58hHxDaJaGXGY3nuvUYFxMzQGbnrxZcFiF6UWMPUsSMy21B6J2Ct8O8EmrFByMxFUN1O
JsJzcpEb8IMP+PeN0RDBe+dIL3ZpbgTqHZruvFFTdHGEcpBNDdDiJ4AvmOfJruRYVKcoYr5j8/y8
jG2he8dAyjSJ5Z15lFtf8Gl1i+XqKb34Y4A/PzVawIxV1IONLWzrAghZRHmgLhCvl1XXXLTsAcMn
Y/aCNK/aYoILcF+6G3UTcAzl5ypOIxZY1tYhzYjuB2OTyj342QMXdEl1k1tG1y0lnxs2tO0d5n3u
IYDCVqPzs0TzuFKMYcoEnKCYmGI14aN69RDqVdsw8ldkngnkZaKmBX4ukfZ+C5dKELX0H0t5QJpY
UGwpMBKdroD8L3aoHa0wgWvPFRChkTvUO2MdYiiM8ppkr0mqJEoLpcVscxAWrD27e0F7VO2poI8q
qBpXlb3mFNN5jMzKWLwoTR7CXXYNv8kZutWTtjtZF/ADjxZRmVbTR2zsawwZCJQyzEAdOyu5Z8Ep
VgG2vT9FUvSZejABxzHjjubZB3rO442K0rGJgo4S2yOkq5oQPL3mqIWkMwtVgUhZGJ7Wg5nN9Jyw
K+OY8sbmOhsIZfZ90bng4UNqkeX0BsJy3eZsVEn4kOjDyQKRksjOmnOk7zheB4NC+pFhvSry3YRK
DNJHUWmoHPdDEyajQjgdDevofIOyfelTbQCr606YoxQKD09TY0LHXzqSU50pcuDQqCLm75eCg8BS
JS8LlmhTfnsX1CME4hILLB1H0GRwjsIKM5+o+XaCsXtUNwXqzTVQWeWlFXiCFUQZI0Bp3IkrU/XS
15SLpIJxVot2FzY8g7jXaTtvJfHLLcHGXYqZUywSmyc/ZpTMrPu+YEVLq2k319qQPG2GdA2vrd84
32f+LUyz8F5+HfPVAo4tXUtud6L8vXpC0c5/fZ6Hk0AfjAnCof5XTUuSyogJFwRVs3Bzg18L6vlx
V67osxHSnRgRax/KBFwlo2ML5VtAAFS2yMlZmYieEXn+KfZd4UuzF5Ozve8Mq0m9UkVki7pAD53T
UVMISC5uJ8dCm6PbIoqhPKh9jLWljOd5pTRI+ZomuEkpk0BLsb0LDgDPGlIq7NuTE5N0NbxDfJ5m
gJd37yPAPRiKjBtgZ0idE3yM3nvmYhm572Juw9QSxF6u+b9ZK1ErGsMzLrb3jw/mQW+mlzrf+km0
ZaW/nIOf5UJy3ltzlpLqw/v6WbKKxOR7PBC+xloyv13VD5qyYqLUoHdQ21O+gaikZph+jXJrXpkl
4EX/AbAugsbAk25Fm/RYcYffy+WzyM1ZDFh+6/Sc0OWy5ESygqT9hwBUQXdTm2wD27x+fGNYl+sr
suxrPrvAzO7H74za3tfNihA6wwF+Qd4dr1deeegJ6UMJTBKFkuiiBf1TZPfxmYbrhm0eKsmejxJD
VqxchD9m1dVr2I4PQfDhKZdf5olaHnNhoU7ReDWR9IwcyTHLMhahr0h9i3V7U5lBqhAgy6mKNgqI
PQgBGlB6tYSF5sUGM03aXT6sTJq5wGxoh5qtpjKVJSjs1c/ZCg==
`protect end_protected
